module am(IZZ,IAA,IAB,IAC,IAD,IAE,IAF,IAG,IAH,IAI,IAJ,IAK,IAL,IAM,IAN,IAO,IAP,IBA,IBB,IBC,IBD,IBE,IBF,IBG,IBH,IBI,IBJ,IBK,IBL,IBM,IBN,IBO,IBP,ICA,ICB,ICC,ICD,ICE,ICF,ICG,ICH,ICI,ICJ,ICK,ICL,ICM,ICN,ICO,ICP,IDA,IDB,IDC,IDD,IDE,IDF,IDG,IDH,IDI,IDJ,IDK,IDL,IDM,IDN,IDO,IDP,IEA,IEB,IEC,IED,IEE,IEF,IFA,IFB,IFC,IFD,IFE,IFF,IFG,IGA,IGB,IGC,IGD,IGE,IGF,IHA,OAA,OAB,OAC,OAD,OAE,OAF,OAG,OAH,OAI,OAJ,OAK,OAL,OAM,OAN,OAO,OAP,OBA,OBB,OBC,OBD,OBE,OBF,OBG,OBH,OBI,OBJ,OBK,OBL,OBM,OBN,OBO,OBP,OEA,OEB,OEC,OED,OEE,OEF,OFA,OFB,OFC,OFD,OFE,OFF,OGA,OGB,OGC,OGD,OGE,OGF,OHA,OHB,OHC,OHD,OHE,OHF,OIA,OIB,OIC,OID,OIE,OIF,OIG,OIH,OIJ,OIK,OIL,OIM,OJA,OJB,OJC,OJD,OJE,OJF,OJG,OJH,OJI,OJJ,OJK,OJL,OJM,OKA,OKB,OKC,OKD,OKE,OKF,OKG,OKH,OKI,OKJ,OKK,OKL,OKM,OLA,OLB,OLC,OLD,OLE,OLF,OLG,OLH,OLI,OLJ,OLK,OLL,OLM,OMA,OMB,OMC,OMD,OME,OMF,OMG,OMH,OMI,OMJ,OMK,OML,ONA,ONB,ONC,OND,ONE,ONF,ONG,ONH,ONI,ONJ,ONK,ONL,ONM,OOA,OOB,OOC,OOD,OOE,OOF,OOG,OOH,OOI,OOJ,OOK,OOL,OOM,OPA,OPB,OPC,OPD,OPE,OPF,OPG,OPH,OPI,OPJ,OPK,OPL,OPM); 
	// MODULE NAME: AM
	// DESCRIPTION: Address Multiply
	//
	input IZZ,IAA,IAB,IAC,IAD,IAE,IAF,IAG,IAH,IAI,IAJ,IAK,IAL,IAM,IAN,IAO,IAP,IBA,IBB,IBC,IBD,IBE,IBF,IBG,IBH,IBI,IBJ,IBK,IBL,IBM,IBN,IBO,IBP,ICA,ICB,ICC,ICD,ICE,ICF,ICG,ICH,ICI,ICJ,ICK,ICL,ICM,ICN,ICO,ICP,IDA,IDB,IDC,IDD,IDE,IDF,IDG,IDH,IDI,IDJ,IDK,IDL,IDM,IDN,IDO,IDP,IEA,IEB,IEC,IED,IEE,IEF,IFA,IFB,IFC,IFD,IFE,IFF,IFG,IGA,IGB,IGC,IGD,IGE,IGF,IHA; 
	output OAA,OAB,OAC,OAD,OAE,OAF,OAG,OAH,OAI,OAJ,OAK,OAL,OAM,OAN,OAO,OAP,OBA,OBB,OBC,OBD,OBE,OBF,OBG,OBH,OBI,OBJ,OBK,OBL,OBM,OBN,OBO,OBP,OEA,OEB,OEC,OED,OEE,OEF,OFA,OFB,OFC,OFD,OFE,OFF,OGA,OGB,OGC,OGD,OGE,OGF,OHA,OHB,OHC,OHD,OHE,OHF,OIA,OIB,OIC,OID,OIE,OIF,OIG,OIH,OIJ,OIK,OIL,OIM,OJA,OJB,OJC,OJD,OJE,OJF,OJG,OJH,OJI,OJJ,OJK,OJL,OJM,OKA,OKB,OKC,OKD,OKE,OKF,OKG,OKH,OKI,OKJ,OKK,OKL,OKM,OLA,OLB,OLC,OLD,OLE,OLF,OLG,OLH,OLI,OLJ,OLK,OLL,OLM,OMA,OMB,OMC,OMD,OME,OMF,OMG,OMH,OMI,OMJ,OMK,OML,ONA,ONB,ONC,OND,ONE,ONF,ONG,ONH,ONI,ONJ,ONK,ONL,ONM,OOA,OOB,OOC,OOD,OOE,OOF,OOG,OOH,OOI,OOJ,OOK,OOL,OOM,OPA,OPB,OPC,OPD,OPE,OPF,OPG,OPH,OPI,OPJ,OPK,OPL,OPM; 

	reg AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL,AAM,AAN,AAO,AAP,AAQ,ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL,ABM,ABN,ABO,ABP,ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL,ACM,ACN,ACO,ACP,ACQ,ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL,ADM,ADN,ADO,ADP,BAA,BAB,BAC,BAD,BAE,BAF,BAG,BAH,BAI,BAJ,BAK,BAL,BAM,BAN,BAO,BAP,BBA,BBB,BBC,BBD,BBE,BBF,BBG,BBH,BBI,BBJ,BBK,BBL,BBM,BBN,BBO,BBP,DGA,DGC,DGD,dge,DGF,DGG,dgh,DGJ,dgk,DHA,dhb,DHC,dhd,DHE,DHF,DIA,dib,DIC,did,DIE,dif,DIG,DJA,djb,DJC,djd,DJE,djf,DJG,djh,DKA,dkb,DKC,dkd,DKE,dkf,DKG,dkh,DKI,DKJ,DLA,dlb,DLC,dld,DLE,dlf,DLG,dlh,DLI,dlj,DLK,DMA,dmb,DMC,dmd,DME,dmf,DMG,dmh,DMI,dmj,DMK,dml,DNA,dnb,DNC,dnd,DNE,dnf,DNG,dnh,DNI,dnj,DNK,dnl,DNM,DNO,DOA,dob,DOC,dod,DOE,dof,DOG,doh,DOI,doj,DOK,dol,DOM,don,DOO,DPA,dpb,DPC,dpd,DPE,dpf,DPG,dph,DPI,dpj,DPK,dpl,DPM,dpn,DPO,dpp,DQA,dqb,DQC,dqd,DQE,dqf,DQG,dqh,DQI,dqj,DQK,dql,DQM,dqn,DQO,dqp,DQQ,DQR,DRA,drb,DRC,drd,DRE,drf,DRG,drh,DRI,drj,DRK,drl,DRM,drn,DRO,drp,DRQ,drr,DRS,DSA,dsb,DSC,dsd,DSE,dsf,DSG,dsh,DSI,dsj,DSK,dsl,DSM,dsn,DSO,dsp,DSQ,dsr,DSS,dst,DTA,dtb,DTC,dtd,DTE,dtf,DTG,dth,DTI,dtj,DTK,dtl,DTM,dtn,DTO,dtp,DTQ,dtr,DTS,dtt,DTU,DTV,GAA,gab,GAC,gad,GAE,GAF,GBA,gbb,GBC,gbd,GBE,GCA,gcb,GCC,gcd,GCE,GDA,gdb,GDC,gdd,GDE,GEA,geb,GEC,ged,GFA,gfb,GFC,gfd,GFE,GGA,ggb,GGC,ggd,GHA,ghb,GHC,ghd,GHE,GIA,gib,GIC,gid,GJA,gjb,GJC,GJD,GKA,gkb,GKC,gkd,GLA,glb,GLC,GLD,GMA,gmb,GMC,GMD,GNA,gnb,GNC,GND,GOA,gob,GOC,GPA,gpb,GPC,GQA,gqb,GQC,GRA,grb,GRC,GSA,gsb,GSC,GTA,gtb,GUA,gub,GVA,gvb,GWA,GWB,GXA,gxb,GYA,GYB,GZA,GZB,GZD,GZE,GZF,GZH,GZK,GZL,GZM,GZN,JAA,jab,JAC,JBA,jbb,JBC,JCA,jcb,JCC,JDA,jdb,JEA,jeb,JEC,JFA,jfb,JGA,jgb,JGC,JHA,jhb,JIA,jib,JJA,jjb,JKA,jkb,JLA,jlb,JMA,jmb,JNA,JNB,JOA,JOB,JPA,JPB,JQA,JQB,JRA,JRB,JSA,JSB,JTA,JTB,JUA,JUB,JVA,JVB,JWA,JWB,JXA,JXB,JYA,JYB,JZA,JZC,JZD,JZE,JZG,JZI,JZK,JZL,KBA,kbb,KBC,KCA,kcb,KCC,KDA,kdb,KDC,KEA,keb,KFA,kfb,KFC,KGA,kgb,KHA,khb,KHC,KIA,kib,KJA,kjb,KKA,kkb,KLA,klb,KMA,kmb,KNA,knb,KOA,KOB,KPA,KPB,KQA,KQB,KRA,KRB,KSA,KSB,KTA,KTB,KUA,KUB,KVA,KVB,KWA,KWB,KXA,KXB,KYA,KYB,KZA,KZB,KZC,KZE,KZF,KZG,KZI,KZJ,KZL,KZM,MAA,MAB,MAC,MAD,MAE,MAF,MAG,MAH,MAI,MAJ,MAK,MAL,MAM,MAN,MAO,MAP,MBA,MBB,MBC,MBD,MBE,MBF,MBG,MBH,MBI,MBJ,MBK,MBL,MBM,MBN,MBO,MBP,mca,mcb,mcc,mcd,mce,mcf,mcg,mch,mci,mcj,mck,mcl,mcm,mcn,mco,mcp,mda,mdb,mdc,mdd,mde,mdf,mdg,mdh,mdi,MDJ,MDK,MDL,MDM,MDN,MDQ,MEA,MEB,MEC,MED,MEE,MEF,MEH,NAA,NAB,NAC,NAD,NAE,NAF,NAG,NAH,NAI,NAJ,NAK,NAL,NAM,NAN,NAO,NAP,NBA,NBB,NBC,NBD,NBE,NBF,NBG,NBH,NBI,NBJ,NBK,NBL,NBM,NBN,NBO,NBP,NBQ,NEA,NEB,NEC,NED,nee,nef,neg,NEH,nei,nej,nek,nel,nem,nen,neo,nep,nfa,nfb,nfc,nfd,nfe,nff,nfg,nfh,nfi,nfj,nfk,nfl,nfm,nfn,nfo,nfp,OAA,OAB,OAC,OAD,OAE,OAF,OAG,OAH,OAI,OAJ,OAK,OAL,OAM,OAN,OAO,OAP,OBA,OBB,OBC,OBD,OBE,OBF,OBG,OBH,OBI,OBJ,OBK,OBL,OBM,OBN,OBO,OBP,OEA,OEB,OEC,OED,OEE,OEF,OFA,OFB,OFC,OFD,OFE,OFF,oga,ogb,ogc,ogd,oge,ogf,oha,ohb,ohc,ohd,ohe,ohf,oia,oib,oic,oid,oie,oif,oig,oih,oii,oij,oik,oil,oim,OJA,OJB,OJC,OJD,OJE,OJF,OJG,OJH,OJI,OJJ,OJK,OJL,OJM,oka,okb,okc,okd,oke,okf,okg,okh,oki,okj,okk,okl,okm,OLA,OLB,OLC,OLD,OLE,OLF,OLG,OLH,OLI,OLJ,OLK,OLL,OLM,oma,omb,omc,omd,ome,omf,omg,omh,omi,omj,omk,oml,omm,ONA,ONB,ONC,OND,ONE,ONF,ONG,ONH,ONI,ONJ,ONK,ONL,ONM,ooa,oob,ooc,ood,ooe,oof,oog,ooh,ooi,ooj,ook,ool,oom,OPA,OPB,OPC,OPD,OPE,OPF,OPG,OPH,OPI,OPJ,OPK,OPL,OPM,PAB,PAC,PAD,PAE,PAF,PAG,PAH,pai,pak,PAL,PBA,PBB,PBC,PBD,PBE,PBF,PBG,PBH,PBI,PBJ,PBK,PBL,PBM,PBN,PBO,PBP,PCA,PCB,PCC,PCD,PCE,PCF,PCG,PCH,PCI,PCJ,PCK,PCL,PCM,PCN,PCO,PCP,PDE,PDF,PDG,PDH,PDI,PDJ,PDK,PDL,PDM,PDN,PDO,PDP,PEA,PEB,PEC,PED,PEE,PEF,PEG,PEH,PEI,PEJ,PEK,PEL,PEM,PEN,PEO,PEP,PFA,PFB,PFC,PFD,PFE,PFF,PFG,PFH,PFI,PFJ,PFK,PFL,PFM,PFN,PFO,PFP,PGA,PGB,PGC,PGD,PGE,PGF,PGG,PGH,PGI,PGJ,PGK,PGL,PGM,PGN,PGO,PGP,QAA,QAB,QAC,QAD,QAE,QAF,QAG,QAH,QAI,QAJ,QAK,TFA,TFB,TFC,TFD;
	wire CAA,CAB,CAC,CAD,CAE,CAF,CAG,CAH,CAI,CAJ,CAK,CAL,CAM,CAN,CAO,CAP,CBA,CBB,CBC,CBD,CBE,CBF,CBG,CBH,CBI,CBJ,CBK,CBL,CBM,CBN,CBO,CBP,CCA,CCB,CCC,CCD,CCE,CCF,CCG,CCH,CCI,CCJ,CCK,CCL,CCM,CCN,CCO,CDA,CDB,CDC,CDD,CDE,CDF,CDG,CDH,CDI,CDJ,CDK,CDL,CDM,CDN,CDO,CEA,CEB,CEC,CED,CEE,CEF,CEG,CEH,CEI,CEJ,CEK,CEL,CEM,CEN,CFA,CFB,CFC,CFD,CFE,CFF,CFG,CFH,CFI,CFJ,CFK,CFL,CFM,CFN,CGA,CGB,CGC,CGD,CGE,CGF,CGG,CGH,CGI,CGJ,CGK,CGL,CGM,CHA,CHB,CHC,CHD,CHE,CHF,CHG,CHH,CHI,CHJ,CHK,CHL,CHM,CIA,CIB,CIC,CID,CIE,CIF,CIG,CIH,CII,CIJ,CIK,CIL,CJA,CJB,CJC,CJD,CJE,CJF,CJG,CJH,CJI,CJJ,CJK,CJL,CKA,CKB,CKC,CKD,CKE,CKF,CKG,CKH,CKI,CKJ,CKK,CLA,CLB,CLC,CLD,CLE,CLF,CLG,CLH,CLI,CLJ,CLK,CMA,CMB,CMC,CMD,CME,CMF,CMG,CMH,CMI,CMJ,CNA,CNB,CNC,CND,CNE,CNF,CNG,CNH,CNI,CNJ,COA,COB,COC,COD,COE,COF,COG,COH,COI,CPA,CPB,CPC,CPD,CPE,CPF,CPG,CPH,CPI,CQA,CQB,CQC,CQD,CQE,CQF,CQG,CQH,CRA,CRB,CRC,CRD,CRE,CRF,CRG,CRH,CSA,CSB,CSC,CSD,CSE,CSF,CSG,CTA,CTB,CTC,CTD,CTE,CTF,CTG,CUA,CUB,CUC,CUD,CUE,CUF,CVA,CVB,CVC,CVD,CVE,CVF,CWA,CWB,CWC,CWD,CWE,CXA,CXB,CXC,CXD,CXE,CYA,CYB,CYC,CYD,CZA,CZB,CZC,CZD,DAA,DAB,DAC,DBA,DBB,DBC,DCA,DCB,DDA,DDB,DEA,DFA,ECA,ECB,EEA,EEB,EFA,EFB,EGA,egb,EHA,ehb,EIA,eib,EJA,ejb,EKA,ekb,ELA,elb,EMA,emb,EMC,EMD,ENA,enb,ENC,END,EOA,eob,EOC,eod,EPA,epb,EPC,EPD,EQA,eqb,EQC,eqd,ERA,erb,ERC,erd,ESA,esb,ESC,esd,ETA,etb,ETC,etd,EUA,eub,EUC,eud,EUE,EUF,EVA,evb,EVC,evd,EWA,ewb,EWC,ewd,EWE,EWF,EXA,exb,EXC,exd,EXE,EXF,EYA,eyb,EYC,eyd,EYE,eyf,FAA,fab,FAC,fad,FAE,faf,FBA,fbb,FBC,fbd,FBE,fbf,FCA,fcb,FCC,fcd,FCE,fcf,FDA,fdb,FDC,fdd,FDE,fdf,FEA,feb,FEC,fed,FEE,fef,FFA,ffb,FFC,ffd,FFE,fff,FFG,FFH,FGA,fgb,FGC,fgd,FGE,fgf,FGG,FGH,HAA,hab,HAC,HAD,HBA,hbb,HBC,HBD,HCA,hcb,HCD,HCE,HDA,hdb,HDC,HDD,HEA,heb,HFA,hfb,HFC,HFD,HGA,hgb,HHA,hhb,HHC,HHD,HIA,hib,HJA,hjb,HKA,hkb,HLA,hlb,HMA,hmb,HNA,hnb,HOA,hob,HPA,hpb,HQA,hqb,HRA,hrb,HSA,hsb,HTA,HTB,HUA,HUB,HVA,HVB,HWA,HWB,HXA,HXB,HYA,HYB,HZA,HZB,HZE,HZF,LBA,lbb,LBC,lbd,LCA,lcb,LCC,lcd,LDA,LDB,LDC,ldd,LEA,leb,LEC,LED,LFA,lfb,LFC,LFD,LGA,lgb,LGC,LGD,LHA,lhb,LHC,LHD,LIA,lib,LIC,LJA,ljb,LKA,lkb,LLA,llb,LMA,lmb,LNA,lnb,LOA,lob,LPA,lpb,LQA,lqb,LRA,lrb,LSA,lsb,LTA,ltb,LUA,lub,LVA,lvb,LWA,lwb,LXA,lxb,LYA,LYB,LZA,lzb,LZD,lze,LZF,LZG,LZH,LZI,LZJ,LZK,LZL,LZM,LZN,LZO,NHC,NHD,NHE,NIC,NID,NIE,NJC,NJD,NJE,NKC,NKD,NKE,NLC,NLD,NLE,NMC,NMD,NME,NNC,NND,NNE,NPC,NPD,NQC,NQD,NRC,NRD,NSC,NSD,NTC,NTD,NUC,NUD,NVC,NVD,nxb,nxc,nxd,nxe,nxf,nxg,nxi,nxj,nxk,nxl,PAM,ZZI,ZZO;

	assign ZZI = 1'b1;
	assign ZZO = 1'b0;
	assign FGA = ~dtb & dtd & dtf | dtb & ~dtd & dtf | dtb & dtd & ~dtf | ~dtb & ~dtd & ~dtf; 
	assign fgb = ~dtb & dtd & dtf | dtb & ~dtd & dtf | dtb & dtd & ~dtf | dtb & dtd & dtf; 
	assign FGC = ~dth & dtj & dtl | dth & ~dtj & dtl | dth & dtj & ~dtl | ~dth & ~dtj & ~dtl; 
	assign fgd = ~dth & dtj & dtl | dth & ~dtj & dtl | dth & dtj & ~dtl | dth & dtj & dtl; 
	assign FGE = ~dtn & dtp & dtr | dtn & ~dtp & dtr | dtn & dtp & ~dtr | ~dtn & ~dtp & ~dtr; 
	assign fgf = ~dtn & dtp & dtr | dtn & ~dtp & dtr | dtn & dtp & ~dtr | dtn & dtp & dtr; 
	assign FFA = DTA & ~DTC & ~DTE | ~DTA & DTC & ~DTE | ~DTA & ~DTC & DTE | DTA & DTC & DTE; 
	assign ffb = DTA & ~DTC & ~DTE | ~DTA & DTC & ~DTE | ~DTA & ~DTC & DTE | ~DTA & ~DTC & ~DTE; 
	assign FFC = DTG & ~DTI & ~DTK | ~DTG & DTI & ~DTK | ~DTG & ~DTI & DTK | DTG & DTI & DTK; 
	assign ffd = DTG & ~DTI & ~DTK | ~DTG & DTI & ~DTK | ~DTG & ~DTI & DTK | ~DTG & ~DTI & ~DTK; 
	assign FFE = DTM & ~DTO & ~DTQ | ~DTM & DTO & ~DTQ | ~DTM & ~DTO & DTQ | DTM & DTO & DTQ; 
	assign fff = DTM & ~DTO & ~DTQ | ~DTM & DTO & ~DTQ | ~DTM & ~DTO & DTQ | ~DTM & ~DTO & ~DTQ; 
	assign FEA = ~dsb & dsd & dsf | dsb & ~dsd & dsf | dsb & dsd & ~dsf | ~dsb & ~dsd & ~dsf; 
	assign feb = ~dsb & dsd & dsf | dsb & ~dsd & dsf | dsb & dsd & ~dsf | dsb & dsd & dsf; 
	assign FEC = ~dsh & dsj & dsl | dsh & ~dsj & dsl | dsh & dsj & ~dsl | ~dsh & ~dsj & ~dsl; 
	assign fed = ~dsh & dsj & dsl | dsh & ~dsj & dsl | dsh & dsj & ~dsl | dsh & dsj & dsl; 
	assign FEE = ~dsn & dsp & dsr | dsn & ~dsp & dsr | dsn & dsp & ~dsr | ~dsn & ~dsp & ~dsr; 
	assign fef = ~dsn & dsp & dsr | dsn & ~dsp & dsr | dsn & dsp & ~dsr | dsn & dsp & dsr; 
	assign FDA = DSA & ~DSC & ~DSE | ~DSA & DSC & ~DSE | ~DSA & ~DSC & DSE | DSA & DSC & DSE; 
	assign fdb = DSA & ~DSC & ~DSE | ~DSA & DSC & ~DSE | ~DSA & ~DSC & DSE | ~DSA & ~DSC & ~DSE; 
	assign FDC = DSG & ~DSI & ~DSK | ~DSG & DSI & ~DSK | ~DSG & ~DSI & DSK | DSG & DSI & DSK; 
	assign fdd = DSG & ~DSI & ~DSK | ~DSG & DSI & ~DSK | ~DSG & ~DSI & DSK | ~DSG & ~DSI & ~DSK; 
	assign FDE = DSM & ~DSO & ~DSQ | ~DSM & DSO & ~DSQ | ~DSM & ~DSO & DSQ | DSM & DSO & DSQ; 
	assign fdf = DSM & ~DSO & ~DSQ | ~DSM & DSO & ~DSQ | ~DSM & ~DSO & DSQ | ~DSM & ~DSO & ~DSQ; 
	assign FCA = ~drb & drd & drf | drb & ~drd & drf | drb & drd & ~drf | ~drb & ~drd & ~drf; 
	assign fcb = ~drb & drd & drf | drb & ~drd & drf | drb & drd & ~drf | drb & drd & drf; 
	assign FCC = ~drh & drj & drl | drh & ~drj & drl | drh & drj & ~drl | ~drh & ~drj & ~drl; 
	assign fcd = ~drh & drj & drl | drh & ~drj & drl | drh & drj & ~drl | drh & drj & drl; 
	assign FCE = ~drn & drp & drr | drn & ~drp & drr | drn & drp & ~drr | ~drn & ~drp & ~drr; 
	assign fcf = ~drn & drp & drr | drn & ~drp & drr | drn & drp & ~drr | drn & drp & drr; 
	assign FBA = DRA & ~DRC & ~DRE | ~DRA & DRC & ~DRE | ~DRA & ~DRC & DRE | DRA & DRC & DRE; 
	assign fbb = DRA & ~DRC & ~DRE | ~DRA & DRC & ~DRE | ~DRA & ~DRC & DRE | ~DRA & ~DRC & ~DRE; 
	assign CAA = BAA & ACA; 
	assign CAB = BAA & ACC; 
	assign CAC = BAA & ACE; 
	assign CPB = BAP & ACB; 
	assign CPC = BAP & ACD; 
	assign CPD = BAP & ACF; 
	assign CAD = BAA & ACG; 
	assign CAE = BAA & ACI; 
	assign CAF = BAA & ACK; 
	assign CPE = BAP & ACH; 
	assign CPF = BAP & ACJ; 
	assign CPG = BAP & ACL; 
	assign CAG = BAA & ACM; 
	assign CAH = BAA & ACO; 
	assign CAI = BAA & ADA; 
	assign CPH = BAP & ACN; 
	assign CPI = BAP & ACP; 
	assign CQA = BBA & ACA; 
	assign CAJ = BAA & ADC; 
	assign CAK = BAA & ADE; 
	assign CAL = BAA & ADG; 
	assign CQB = BBA & ACC; 
	assign CQC = BBA & ACE; 
	assign CQD = BBA & ACG; 
	assign CAM = BAA & ADI; 
	assign CAN = BAA & ADK; 
	assign CAO = BAA & ADM; 
	assign CQE = BBA & ACI; 
	assign CQF = BBA & ACK; 
	assign CQG = BBA & ACM; 
	assign CAP = BAA & ADO; 
	assign CBA = BAB & ACQ; 
	assign CBB = BAB & ACB; 
	assign CQH = BBA & ACO; 
	assign CRA = BBB & ACQ; 
	assign CRB = BBB & ACB; 
	assign CBC = BAB & ACD; 
	assign CBD = BAB & ACF; 
	assign CBE = BAB & ACH; 
	assign CRC = BBB & ACD; 
	assign CRD = BBB & ACF; 
	assign CRE = BBB & ACH; 
	assign CBF = BAB & ACJ; 
	assign CBG = BAB & ACL; 
	assign CBH = BAB & ACN; 
	assign CRF = BBB & ACJ; 
	assign CRG = BBB & ACL; 
	assign CRH = BBB & ACN; 
	assign EPD = ~dlh & ~dlj; 
	assign END = ~dkh & DKJ; 
	assign FFG = DTS & ~DTU | ~DTS & DTU; 
	assign FGG = ~dtt & ~DTV | dtt & DTV; 
	assign EUF = DOM & DOO; 
	assign EXF = ~dpn & ~dpp; 
	assign FGH = ~dtt & DTV; 
	assign EWF = DPO & DPM ; 
	assign ECA = DGD & ~DGF | ~DGD & DGF; 
	assign EEA = DGG & ~DGJ | ~DGG & DGJ; 
	assign EMC = DKG & ~DKI | ~DKG & DKI; 
	assign EPC = ~dlh & dlj | dlh & ~dlj; 
	assign EXE = ~dpn & dpp | dpn & ~dpp; 
	assign FBC = DRG & ~DRI & ~DRK | ~DRG & DRI & ~DRK | ~DRG & ~DRI & DRK | DRG & DRI & DRK; 
	assign fbd = DRG & ~DRI & ~DRK | ~DRG & DRI & ~DRK | ~DRG & ~DRI & DRK | ~DRG & ~DRI & ~DRK; 
	assign FBE = DRM & ~DRO & ~DRQ | ~DRM & DRO & ~DRQ | ~DRM & ~DRO & DRQ | DRM & DRO & DRQ; 
	assign fbf = DRM & ~DRO & ~DRQ | ~DRM & DRO & ~DRQ | ~DRM & ~DRO & DRQ | ~DRM & ~DRO & ~DRQ; 
	assign FAA = ~dqb & dqd & dqf | dqb & ~dqd & dqf | dqb & dqd & ~dqf | ~dqb & ~dqd & ~dqf; 
	assign fab = ~dqb & dqd & dqf | dqb & ~dqd & dqf | dqb & dqd & ~dqf | dqb & dqd & dqf; 
	assign FAC = ~dqh & dqj & dql | dqh & ~dqj & dql | dqh & dqj & ~dql | ~dqh & ~dqj & ~dql; 
	assign fad = ~dqh & dqj & dql | dqh & ~dqj & dql | dqh & dqj & ~dql | dqh & dqj & dql; 
	assign FAE = ~dqn & dqp & ~DQR | dqn & ~dqp & ~DQR | dqn & dqp & DQR | ~dqn & ~dqp & DQR; 
	assign faf = ~dqn & dqp & ~DQR | dqn & ~dqp & ~DQR | dqn & dqp & DQR | dqn & dqp & ~DQR; 
	assign EYA = DQA & ~DQC & ~DQE | ~DQA & DQC & ~DQE | ~DQA & ~DQC & DQE | DQA & DQC & DQE; 
	assign eyb = DQA & ~DQC & ~DQE | ~DQA & DQC & ~DQE | ~DQA & ~DQC & DQE | ~DQA & ~DQC & ~DQE; 
	assign HAC = ~gbb & gbd | gbb & ~gbd; 
	assign EYC = DQG & ~DQI & ~DQK | ~DQG & DQI & ~DQK | ~DQG & ~DQI & DQK | DQG & DQI & DQK; 
	assign eyd = DQG & ~DQI & ~DQK | ~DQG & DQI & ~DQK | ~DQG & ~DQI & DQK | ~DQG & ~DQI & ~DQK; 
	assign EYE = DQM & ~DQO & ~DQQ | ~DQM & DQO & ~DQQ | ~DQM & ~DQO & DQQ | DQM & DQO & DQQ; 
	assign eyf = DQM & ~DQO & ~DQQ | ~DQM & DQO & ~DQQ | ~DQM & ~DQO & DQQ | ~DQM & ~DQO & ~DQQ; 
	assign HBC = ~gcb & gcd | gcb & ~gcd; 
	assign EXA = ~dpb & dpd & dpf | dpb & ~dpd & dpf | dpb & dpd & ~dpf | ~dpb & ~dpd & ~dpf; 
	assign exb = ~dpb & dpd & dpf | dpb & ~dpd & dpf | dpb & dpd & ~dpf | dpb & dpd & dpf; 
	assign EXC = ~dph & dpj & dpl | dph & ~dpj & dpl | dph & dpj & ~dpl | ~dph & ~dpj & ~dpl; 
	assign exd = ~dph & dpj & dpl | dph & ~dpj & dpl | dph & dpj & ~dpl | dph & dpj & dpl; 
	assign HCD = ~gdb & gdd | gdb & ~gdd; 
	assign EWA = DPA & ~DPC & ~DPE | ~DPA & DPC & ~DPE | ~DPA & ~DPC & DPE | DPA & DPC & DPE; 
	assign ewb = DPA & ~DPC & ~DPE | ~DPA & DPC & ~DPE | ~DPA & ~DPC & DPE | ~DPA & ~DPC & ~DPE; 
	assign EWC = DPG & ~DPI & ~DPK | ~DPG & DPI & ~DPK | ~DPG & ~DPI & DPK | DPG & DPI & DPK; 
	assign ewd = DPG & ~DPI & ~DPK | ~DPG & DPI & ~DPK | ~DPG & ~DPI & DPK | ~DPG & ~DPI & ~DPK; 
	assign EWE = DPM & ~DPO | ~DPM & DPO; 
	assign EVA = ~dob & dod & dof | dob & ~dod & dof | dob & dod & ~dof | ~dob & ~dod & ~dof; 
	assign evb = ~dob & dod & dof | dob & ~dod & dof | dob & dod & ~dof | dob & dod & dof; 
	assign EVC = ~doh & doj & dol | doh & ~doj & dol | doh & doj & ~dol | ~doh & ~doj & ~dol; 
	assign evd = ~doh & doj & dol | doh & ~doj & dol | doh & doj & ~dol | doh & doj & dol; 
	assign EUA = DOA & ~DOC & ~DOE | ~DOA & DOC & ~DOE | ~DOA & ~DOC & DOE | DOA & DOC & DOE; 
	assign eub = DOA & ~DOC & ~DOE | ~DOA & DOC & ~DOE | ~DOA & ~DOC & DOE | ~DOA & ~DOC & ~DOE; 
	assign CBI = BAB & ACP; 
	assign CBJ = BAB & ADB; 
	assign CBK = BAB & ADD; 
	assign CSA = BBC & ACA; 
	assign CSB = BBC & ACC; 
	assign CSC = BBC & ACE; 
	assign CBL = BAB & ADF; 
	assign CBM = BAB & ADH; 
	assign CBN = BAB & ADJ; 
	assign CSD = BBC & ACG; 
	assign CSE = BBC & ACI; 
	assign CSF = BBC & ACK; 
	assign CBO = BAB & ADL; 
	assign CBP = BAB & ADN; 
	assign CCA = BAC & ACA; 
	assign CSG = BBC & ACM; 
	assign CTA = BBD & ACQ; 
	assign CTB = BBD & ACB; 
	assign CCB = BAC & ACC; 
	assign CCC = BAC & ACE; 
	assign CCD = BAC & ACG; 
	assign CTC = BBD & ACD; 
	assign CTD = BBD & ACF; 
	assign CTE = BBD & ACH; 
	assign CCE = BAC & ACI; 
	assign CCF = BAC & ACK; 
	assign CCG = BAC & ACM; 
	assign CTF = BBD & ACJ; 
	assign CTG = BBD & ACL; 
	assign CUA = BBE & ACA; 
	assign HBD = ~gcb & ~gcd; 
	assign HZF = GZF & GZN; 
	assign HCE = ~gdb & ~gdd; 
	assign CCH = BAC & ACO; 
	assign CCI = BAC & ADA; 
	assign CCJ = BAC & ADC; 
	assign CUB = BBE & ACC; 
	assign CUC = BBE & ACE; 
	assign CUD = BBE & ACG; 
	assign CCK = BAC & ADE; 
	assign CCL = BAC & ADG; 
	assign CCM = BAC & ADI; 
	assign CUE = BBE & ACI; 
	assign CUF = BBE & ACK; 
	assign CVA = BBF & ACQ; 
	assign CCN = BAC & ADK; 
	assign CCO = BAC & ADM; 
	assign CDA = BAD & ACQ; 
	assign CVB = BBF & ACB; 
	assign CVC = BBF & ACD; 
	assign CVD = BBF & ACF; 
	assign LFC = ~kgb & ~KFC | kgb & KFC; 
	assign HDC = ~geb & ged | geb & ~ged; 
	assign HDD = ~ged & ~geb ; 
	assign EUC = DOG & ~DOI & ~DOK | ~DOG & DOI & ~DOK | ~DOG & ~DOI & DOK | DOG & DOI & DOK; 
	assign eud = DOG & ~DOI & ~DOK | ~DOG & DOI & ~DOK | ~DOG & ~DOI & DOK | ~DOG & ~DOI & ~DOK; 
	assign ETA = ~dnb & dnd & dnf | dnb & ~dnd & dnf | dnb & dnd & ~dnf | ~dnb & ~dnd & ~dnf; 
	assign etb = ~dnb & dnd & dnf | dnb & ~dnd & dnf | dnb & dnd & ~dnf | dnb & dnd & dnf; 
	assign ETC = ~dnh & dnj & dnl | dnh & ~dnj & dnl | dnh & dnj & ~dnl | ~dnh & ~dnj & ~dnl; 
	assign etd = ~dnh & dnj & dnl | dnh & ~dnj & dnl | dnh & dnj & ~dnl | dnh & dnj & dnl; 
	assign ESA = DNA & ~DNC & ~DNE | ~DNA & DNC & ~DNE | ~DNA & ~DNC & DNE | DNA & DNC & DNE; 
	assign esb = DNA & ~DNC & ~DNE | ~DNA & DNC & ~DNE | ~DNA & ~DNC & DNE | ~DNA & ~DNC & ~DNE; 
	assign NTD = NBE & NBF & NBG | NBG & ~nff | ~nfg; 
	assign ESC = DNG & ~DNI & ~DNK | ~DNG & DNI & ~DNK | ~DNG & ~DNI & DNK | DNG & DNI & DNK; 
	assign esd = DNG & ~DNI & ~DNK | ~DNG & DNI & ~DNK | ~DNG & ~DNI & DNK | ~DNG & ~DNI & ~DNK; 
	assign ERA = ~dmb & dmd & dmf | dmb & ~dmd & dmf | dmb & dmd & ~dmf | ~dmb & ~dmd & ~dmf; 
	assign erb = ~dmb & dmd & dmf | dmb & ~dmd & dmf | dmb & dmd & ~dmf | dmb & dmd & dmf; 
	assign ERC = ~dmh & dmj & dml | dmh & ~dmj & dml | dmh & dmj & ~dml | ~dmh & ~dmj & ~dml; 
	assign erd = ~dmh & dmj & dml | dmh & ~dmj & dml | dmh & dmj & ~dml | dmh & dmj & dml; 
	assign EQA = DMA & ~DMC & ~DME | ~DMA & DMC & ~DME | ~DMA & ~DMC & DME | DMA & DMC & DME; 
	assign eqb = DMA & ~DMC & ~DME | ~DMA & DMC & ~DME | ~DMA & ~DMC & DME | ~DMA & ~DMC & ~DME; 
	assign HAD = ~gbb & ~gbd; 
	assign EQC = DMG & ~DMI & ~DMK | ~DMG & DMI & ~DMK | ~DMG & ~DMI & DMK | DMG & DMI & DMK; 
	assign eqd = DMG & ~DMI & ~DMK | ~DMG & DMI & ~DMK | ~DMG & ~DMI & DMK | ~DMG & ~DMI & ~DMK; 
	assign EPA = ~dlb & dld & dlf | dlb & ~dld & dlf | dlb & dld & ~dlf | ~dlb & ~dld & ~dlf; 
	assign epb = ~dlb & dld & dlf | dlb & ~dld & dlf | dlb & dld & ~dlf | dlb & dld & dlf; 
	assign EOA = DLA & ~DLC & ~DLE | ~DLA & DLC & ~DLE | ~DLA & ~DLC & DLE | DLA & DLC & DLE; 
	assign eob = DLA & ~DLC & ~DLE | ~DLA & DLC & ~DLE | ~DLA & ~DLC & DLE | ~DLA & ~DLC & ~DLE; 
	assign EOC = DLG & ~DLI & ~DLK | ~DLG & DLI & ~DLK | ~DLG & ~DLI & DLK | DLG & DLI & DLK; 
	assign eod = DLG & ~DLI & ~DLK | ~DLG & DLI & ~DLK | ~DLG & ~DLI & DLK | ~DLG & ~DLI & ~DLK; 
	assign ENA = ~dkb & dkd & dkf | dkb & ~dkd & dkf | dkb & dkd & ~dkf | ~dkb & ~dkd & ~dkf; 
	assign enb = ~dkb & dkd & dkf | dkb & ~dkd & dkf | dkb & dkd & ~dkf | dkb & dkd & dkf; 
	assign EMA = DKA & ~DKC & ~DKE | ~DKA & DKC & ~DKE | ~DKA & ~DKC & DKE | DKA & DKC & DKE; 
	assign emb = DKA & ~DKC & ~DKE | ~DKA & DKC & ~DKE | ~DKA & ~DKC & DKE | ~DKA & ~DKC & ~DKE; 
	assign ELA = ~djb & djd & djf | djb & ~djd & djf | djb & djd & ~djf | ~djb & ~djd & ~djf; 
	assign elb = ~djb & djd & djf | djb & ~djd & djf | djb & djd & ~djf | djb & djd & djf; 
	assign EKA = DJA & ~DJE & ~DJC | ~DJA & DJE & ~DJC | ~DJA & ~DJE & DJC | DJA & DJE & DJC; 
	assign ekb = DJA & ~DJE & ~DJC | ~DJA & DJE & ~DJC | ~DJA & ~DJE & DJC | ~DJA & ~DJE & ~DJC; 
	assign CDB = BAD & ACB; 
	assign CDC = BAD & ACD; 
	assign CDD = BAD & ACF; 
	assign CVE = BBF & ACH; 
	assign CVF = BBF & ACJ; 
	assign CWA = BBG & ACA; 
	assign CDE = BAD & ACH; 
	assign CDF = BAD & ACJ; 
	assign CDG = BAD & ACL; 
	assign CWB = BBG & ACC; 
	assign CWC = BBG & ACE; 
	assign CWD = BBG & ACG; 
	assign CDH = BAD & ACN; 
	assign CDI = BAD & ACP; 
	assign CDJ = BAD & ADB; 
	assign CWE = BBG & ACI; 
	assign CXA = BBH & ACQ; 
	assign CXB = BBH & ACB; 
	assign CDK = BAD & ADD; 
	assign CDL = BAD & ADF; 
	assign CDM = BAD & ADH; 
	assign CXC = BBH & ACD; 
	assign CXD = BBH & ACF; 
	assign CXE = BBH & ACH; 
	assign CDN = BAD & ADJ; 
	assign CDO = BAD & ADL; 
	assign CEA = BAE & ACA; 
	assign CYA = BBI & ACA; 
	assign CYB = BBI & ACC; 
	assign CYC = BBI & ACE; 
	assign CEB = BAE & ACC; 
	assign CEC = BAE & ACE; 
	assign CED = BAE & ACG; 
	assign CYD = BBI & ACG; 
	assign CZA = BBJ & ACQ; 
	assign CZB = BBJ & ACB; 
	assign CEE = BAE & ACI; 
	assign CEF = BAE & ACK; 
	assign CEG = BAE & ACM; 
	assign CZC = BBJ & ACD; 
	assign CZD = BBJ & ACF; 
	assign DAA = BBK & ACA; 
	assign CEH = BAE & ACO; 
	assign CEI = BAE & ADA; 
	assign CEJ = BAE & ADC; 
	assign DAB = BBK & ACC; 
	assign DAC = BBK & ACE; 
	assign DBA = BBL & ACQ; 
	assign HTB = GTA & ~gub; 
	assign PAM = PAL & ~pai; 
	assign HOA = GOA & gpb & ~GOC | ~GOA & ~gpb & ~GOC | ~GOA & gpb & GOC | GOA & ~gpb & GOC; 
	assign hob = GOA & gpb & ~GOC | ~GOA & ~gpb & ~GOC | ~GOA & gpb & GOC | ~GOA & gpb & ~GOC; 
	assign HRA = GRA & gsb & ~GRC | ~GRA & ~gsb & ~GRC | ~GRA & gsb & GRC | GRA & ~gsb & GRC; 
	assign hrb = GRA & gsb & ~GRC | ~GRA & ~gsb & ~GRC | ~GRA & gsb & GRC | ~GRA & gsb & ~GRC; 
	assign HTA = GTA & gub | ~GTA & ~gub; 
	assign HUA = GUA & gvb | ~GUA & ~gvb; 
	assign HUB = GUA & ~gvb; 
	assign HVB = GVA & GWB; 
	assign HWB = GWA & ~gxb; 
	assign HVA = GVA & ~GWB | ~GVA & GWB; 
	assign HWA = GWA & gxb | ~GWA & ~gxb; 
	assign HZA = GZA & ~GZE | ~GZA & GZE; 
	assign HZB = GZA & GZE; 
	assign NQC = NAI & NAJ | ~nej; 
	assign NQD = NAI & NAJ & NAK | NAK & ~nej | ~nek; 
	assign NPD = NAE & NAF & NAG | NAG & ~nef | ~neg; 
	assign NPC = NAE & NAF | ~nef; 
	assign EJA = ~dib & did & dif | dib & ~did & dif | dib & did & ~dif | ~dib & ~did & ~dif; 
	assign ejb = ~dib & did & dif | dib & ~did & dif | dib & did & ~dif | dib & did & dif; 
	assign EIA = DIA & ~DIC & ~DIE | ~DIA & DIC & ~DIE | ~DIA & ~DIC & DIE | DIA & DIC & DIE; 
	assign eib = DIA & ~DIC & ~DIE | ~DIA & DIC & ~DIE | ~DIA & ~DIC & DIE | ~DIA & ~DIC & ~DIE; 
	assign EHA = ~dhb & dhd & ~DHF | dhb & ~dhd & ~DHF | dhb & dhd & DHF | ~dhb & ~dhd & DHF; 
	assign ehb = ~dhb & dhd & ~DHF | dhb & ~dhd & ~DHF | dhb & dhd & DHF | dhb & dhd & ~DHF; 
	assign EGA = DHA & ~DHC & ~DHE | ~DHA & DHC & ~DHE | ~DHA & ~DHC & DHE | DHA & DHC & DHE; 
	assign egb = DHA & ~DHC & ~DHE | ~DHA & DHC & ~DHE | ~DHA & ~DHC & DHE | ~DHA & ~DHC & ~DHE; 
	assign HFC = ~ggb & ggd | ggb & ~ggd; 
	assign HAA = GAA & ~GAC & ~GAE | ~GAA & GAC & ~GAE | ~GAA & ~GAC & GAE | GAA & GAC & GAE; 
	assign hab = GAA & ~GAC & ~GAE | ~GAA & GAC & ~GAE | ~GAA & ~GAC & GAE | ~GAA & ~GAC & ~GAE; 
	assign HBA = GBA & ~GBC & ~GBE | ~GBA & GBC & ~GBE | ~GBA & ~GBC & GBE | GBA & GBC & GBE; 
	assign hbb = GBA & ~GBC & ~GBE | ~GBA & GBC & ~GBE | ~GBA & ~GBC & GBE | ~GBA & ~GBC & ~GBE; 
	assign HFD = ~ggd & ~ggb ; 
	assign HCA = GCA & ~GCC & ~GCE | ~GCA & GCC & ~GCE | ~GCA & ~GCC & GCE | GCA & GCC & GCE; 
	assign hcb = GCA & ~GCC & ~GCE | ~GCA & GCC & ~GCE | ~GCA & ~GCC & GCE | ~GCA & ~GCC & ~GCE; 
	assign HDA = GDA & ~GDC & ~GDE | ~GDA & GDC & ~GDE | ~GDA & ~GDC & GDE | GDA & GDC & GDE; 
	assign hdb = GDA & ~GDC & ~GDE | ~GDA & GDC & ~GDE | ~GDA & ~GDC & GDE | ~GDA & ~GDC & ~GDE; 
	assign HHC = ~gib & gid | gib & ~gid; 
	assign HEA = GEA & ~GEC & gfb | ~GEA & GEC & gfb | ~GEA & ~GEC & ~gfb | GEA & GEC & ~gfb; 
	assign heb = GEA & ~GEC & gfb | ~GEA & GEC & gfb | ~GEA & ~GEC & ~gfb | ~GEA & ~GEC & gfb; 
	assign HFA = GFA & ~GFC & ~GFE | ~GFA & GFC & ~GFE | ~GFA & ~GFC & GFE | GFA & GFC & GFE; 
	assign hfb = GFA & ~GFC & ~GFE | ~GFA & GFC & ~GFE | ~GFA & ~GFC & GFE | ~GFA & ~GFC & ~GFE; 
	assign HHD = ~gid & ~gib ; 
	assign HGA = GGA & ~GGC & ghb | ~GGA & GGC & ghb | ~GGA & ~GGC & ~ghb | GGA & GGC & ~ghb; 
	assign hgb = GGA & ~GGC & ghb | ~GGA & GGC & ghb | ~GGA & ~GGC & ~ghb | ~GGA & ~GGC & ghb; 
	assign HHA = GHA & ~GHC & ~GHE | ~GHA & GHC & ~GHE | ~GHA & ~GHC & GHE | GHA & GHC & GHE; 
	assign hhb = GHA & ~GHC & ~GHE | ~GHA & GHC & ~GHE | ~GHA & ~GHC & GHE | ~GHA & ~GHC & ~GHE; 
	assign HIA = GIA & ~GIC & gjb | ~GIA & GIC & gjb | ~GIA & ~GIC & ~gjb | GIA & GIC & ~gjb; 
	assign hib = GIA & ~GIC & gjb | ~GIA & GIC & gjb | ~GIA & ~GIC & ~gjb | ~GIA & ~GIC & gjb; 
	assign HJA = GJA & ~GJC & gkb | ~GJA & GJC & gkb | ~GJA & ~GJC & ~gkb | GJA & GJC & ~gkb; 
	assign hjb = GJA & ~GJC & gkb | ~GJA & GJC & gkb | ~GJA & ~GJC & ~gkb | ~GJA & ~GJC & gkb; 
	assign HKA = GKA & ~GKC & glb | ~GKA & GKC & glb | ~GKA & ~GKC & ~glb | GKA & GKC & ~glb; 
	assign hkb = GKA & ~GKC & glb | ~GKA & GKC & glb | ~GKA & ~GKC & ~glb | ~GKA & ~GKC & glb; 
	assign HLA = GLA & ~GLC & gmb | ~GLA & GLC & gmb | ~GLA & ~GLC & ~gmb | GLA & GLC & ~gmb; 
	assign hlb = GLA & ~GLC & gmb | ~GLA & GLC & gmb | ~GLA & ~GLC & ~gmb | ~GLA & ~GLC & gmb; 
	assign CEK = BAE & ADE; 
	assign CEL = BAE & ADG; 
	assign CEM = BAE & ADI; 
	assign DBB = BBL & ACB; 
	assign DBC = BBL & ACD; 
	assign DCA = BBM & ACA; 
	assign CEN = BAE & ADK; 
	assign CFA = BAF & ACQ; 
	assign CFB = BAF & ACB; 
	assign DCB = BBM & ACC; 
	assign DDA = BBN & ACQ; 
	assign DDB = BBN & ACB; 
	assign CFC = BAF & ACD; 
	assign CFD = BAF & ACF; 
	assign CFE = BAF & ACH; 
	assign DEA = BBO & ACA; 
	assign DFA = BBP & ACQ; 
	assign CFF = BAF & ACJ; 
	assign CFG = BAF & ACL; 
	assign CFH = BAF & ACN; 
	assign NSC = NBA & NBB | ~nfb; 
	assign NSD = NBA & NBB & NBC | NBC & ~nfb | ~nfc; 
	assign CFI = BAF & ACP; 
	assign CFJ = BAF & ADB; 
	assign CFK = BAF & ADD; 
	assign CFL = BAF & ADF; 
	assign CFM = BAF & ADH; 
	assign CFN = BAF & ADJ; 
	assign nxb = ~NAE | ~NAF | ~NAG | ~NAH;
	assign CGA = BAG & ACA; 
	assign CGB = BAG & ACC; 
	assign CGC = BAG & ACE; 
	assign EFA = ~dgh & dgk | dgh & ~dgk; 
	assign CGD = BAG & ACG; 
	assign CGE = BAG & ACI; 
	assign CGF = BAG & ACK; 
	assign HZE = GZF & ~GZN | ~GZF & GZN; 
	assign nxc = ~NAI | ~NAJ | ~NAK | ~NAL;
	assign nxd = ~NAM | ~NAN | ~NAO | ~NAP;
	assign nxe = ~NBA | ~NBB | ~NBC | ~NBD;
	assign nxf = ~NBE | ~NBF | ~NBG | ~NBH;
	assign NNC = ~nfm & NBN | ~nfn; 
	assign HMA = GMA & ~GMC & gnb | ~GMA & GMC & gnb | ~GMA & ~GMC & ~gnb | GMA & GMC & ~gnb; 
	assign hmb = GMA & ~GMC & gnb | ~GMA & GMC & gnb | ~GMA & ~GMC & ~gnb | ~GMA & ~GMC & gnb; 
	assign HNA = GNA & ~GNC & gob | ~GNA & GNC & gob | ~GNA & ~GNC & ~gob | GNA & GNC & ~gob; 
	assign hnb = GNA & ~GNC & gob | ~GNA & GNC & gob | ~GNA & ~GNC & ~gob | ~GNA & ~GNC & gob; 
	assign HPA = GPA & ~GPC & gqb | ~GPA & GPC & gqb | ~GPA & ~GPC & ~gqb | GPA & GPC & ~gqb; 
	assign hpb = GPA & ~GPC & gqb | ~GPA & GPC & gqb | ~GPA & ~GPC & ~gqb | ~GPA & ~GPC & gqb; 
	assign HQA = GQA & ~GQC & grb | ~GQA & GQC & grb | ~GQA & ~GQC & ~grb | GQA & GQC & ~grb; 
	assign hqb = GQA & ~GQC & grb | ~GQA & GQC & grb | ~GQA & ~GQC & ~grb | ~GQA & ~GQC & grb; 
	assign HSA = GSA & ~GSC & gtb | ~GSA & GSC & gtb | ~GSA & ~GSC & ~gtb | GSA & GSC & ~gtb; 
	assign hsb = GSA & ~GSC & gtb | ~GSA & GSC & gtb | ~GSA & ~GSC & ~gtb | ~GSA & ~GSC & gtb; 
	assign LED = KEA & ~kfb; 
	assign LDB = JDA & ~jeb; 
	assign LBA = JBA & ~JBC & ~KBA | ~JBA & JBC & ~KBA | ~JBA & ~JBC & KBA | JBA & JBC & KBA; 
	assign lbb = JBA & ~JBC & ~KBA | ~JBA & JBC & ~KBA | ~JBA & ~JBC & KBA | ~JBA & ~JBC & ~KBA; 
	assign LBC = KBC & kcb & jcb | ~KBC & ~kcb & jcb | ~KBC & kcb & ~jcb | KBC & ~kcb & ~jcb; 
	assign lbd = KBC & kcb & jcb | ~KBC & ~kcb & jcb | ~KBC & kcb & ~jcb | ~KBC & kcb & jcb; 
	assign LCA = JCA & ~JCC & ~KCA | ~JCA & JCC & ~KCA | ~JCA & ~JCC & KCA | JCA & JCC & KCA; 
	assign lcb = JCA & ~JCC & ~KCA | ~JCA & JCC & ~KCA | ~JCA & ~JCC & KCA | ~JCA & ~JCC & ~KCA; 
	assign LCC = KCA & ~KCC & jdb | ~KCA & KCC & jdb | ~KCA & ~KCC & ~jdb | KCA & KCC & ~jdb; 
	assign lcd = KCA & ~KCC & jdb | ~KCA & KCC & jdb | ~KCA & ~KCC & ~jdb | ~KCA & ~KCC & jdb; 
	assign LDA = JDA & jeb | ~JDA & ~jeb; 
	assign LDC = KDA & ~KDC & keb | ~KDA & KDC & keb | ~KDA & ~KDC & ~keb | KDA & KDC & ~keb; 
	assign ldd = KDA & ~KDC & keb | ~KDA & KDC & keb | ~KDA & ~KDC & ~keb | ~KDA & ~KDC & keb; 
	assign LEA = JEA & ~JEC & jfb | ~JEA & JEC & jfb | ~JEA & ~JEC & ~jfb | JEA & JEC & ~jfb; 
	assign leb = JEA & ~JEC & jfb | ~JEA & JEC & jfb | ~JEA & ~JEC & ~jfb | ~JEA & ~JEC & jfb; 
	assign LEC = KEA & kfb | ~KEA & ~kfb; 
	assign LFA = JFA & jgb & ~KFA | ~JFA & ~jgb & ~KFA | ~JFA & jgb & KFA | JFA & ~jgb & KFA; 
	assign lfb = JFA & jgb & ~KFA | ~JFA & ~jgb & ~KFA | ~JFA & jgb & KFA | ~JFA & jgb & ~KFA; 
	assign LGA = JGA & ~JGC & jhb | ~JGA & JGC & jhb | ~JGA & ~JGC & ~jhb | JGA & JGC & ~jhb; 
	assign lgb = JGA & ~JGC & jhb | ~JGA & JGC & jhb | ~JGA & ~JGC & ~jhb | ~JGA & ~JGC & jhb; 
	assign CGG = BAG & ACM; 
	assign CGH = BAG & ACO; 
	assign CGI = BAG & ADA; 
	assign CGJ = BAG & ADC; 
	assign CGK = BAG & ADE; 
	assign CGL = BAG & ADG; 
	assign CGM = BAG & ADI; 
	assign CHA = BAH & ACQ; 
	assign CHB = BAH & ACB; 
	assign CHC = BAH & ACD; 
	assign CHD = BAH & ACF; 
	assign CHE = BAH & ACH; 
	assign CHF = BAH & ACJ; 
	assign CHG = BAH & ACL; 
	assign CHH = BAH & ACN; 
	assign CHI = BAH & ACP; 
	assign CHJ = BAH & ADB; 
	assign CHK = BAH & ADD; 
	assign CHL = BAH & ADF; 
	assign CHM = BAH & ADH; 
	assign CIA = BAI & ACA; 
	assign CIB = BAI & ACC; 
	assign CIC = BAI & ACE; 
	assign CID = BAI & ACG; 
	assign LGC = KGA & khb | ~KGA & ~khb; 
	assign LHA = JHA & jib & ~KHA | ~JHA & ~jib & ~KHA | ~JHA & jib & KHA | JHA & ~jib & KHA; 
	assign lhb = JHA & jib & ~KHA | ~JHA & ~jib & ~KHA | ~JHA & jib & KHA | ~JHA & jib & ~KHA; 
	assign LIA = JIA & jjb & ~KIA | ~JIA & ~jjb & ~KIA | ~JIA & jjb & KIA | JIA & ~jjb & KIA; 
	assign lib = JIA & jjb & ~KIA | ~JIA & ~jjb & ~KIA | ~JIA & jjb & KIA | ~JIA & jjb & ~KIA; 
	assign LJA = JJA & jkb & ~KJA | ~JJA & ~jkb & ~KJA | ~JJA & jkb & KJA | JJA & ~jkb & KJA; 
	assign ljb = JJA & jkb & ~KJA | ~JJA & ~jkb & ~KJA | ~JJA & jkb & KJA | ~JJA & jkb & ~KJA; 
	assign LKA = JKA & jlb & ~KKA | ~JKA & ~jlb & ~KKA | ~JKA & jlb & KKA | JKA & ~jlb & KKA; 
	assign lkb = JKA & jlb & ~KKA | ~JKA & ~jlb & ~KKA | ~JKA & jlb & KKA | ~JKA & jlb & ~KKA; 
	assign LLA = JLA & jmb & ~KLA | ~JLA & ~jmb & ~KLA | ~JLA & jmb & KLA | JLA & ~jmb & KLA; 
	assign llb = JLA & jmb & ~KLA | ~JLA & ~jmb & ~KLA | ~JLA & jmb & KLA | ~JLA & jmb & ~KLA; 
	assign NTC = NBE & NBF | ~nff; 
	assign LMA = JMA & ~JNB & ~KMA | ~JMA & JNB & ~KMA | ~JMA & ~JNB & KMA | JMA & JNB & KMA; 
	assign lmb = JMA & ~JNB & ~KMA | ~JMA & JNB & ~KMA | ~JMA & ~JNB & KMA | ~JMA & ~JNB & ~KMA; 
	assign LNA = JNA & ~JOB & ~KNA | ~JNA & JOB & ~KNA | ~JNA & ~JOB & KNA | JNA & JOB & KNA; 
	assign lnb = JNA & ~JOB & ~KNA | ~JNA & JOB & ~KNA | ~JNA & ~JOB & KNA | ~JNA & ~JOB & ~KNA; 
	assign LOA = JOA & ~JPB & ~KOA | ~JOA & JPB & ~KOA | ~JOA & ~JPB & KOA | JOA & JPB & KOA; 
	assign lob = JOA & ~JPB & ~KOA | ~JOA & JPB & ~KOA | ~JOA & ~JPB & KOA | ~JOA & ~JPB & ~KOA; 
	assign LPA = JPA & ~JQB & ~KPA | ~JPA & JQB & ~KPA | ~JPA & ~JQB & KPA | JPA & JQB & KPA; 
	assign lpb = JPA & ~JQB & ~KPA | ~JPA & JQB & ~KPA | ~JPA & ~JQB & KPA | ~JPA & ~JQB & ~KPA; 
	assign LQA = JQA & ~JRB & ~KQA | ~JQA & JRB & ~KQA | ~JQA & ~JRB & KQA | JQA & JRB & KQA; 
	assign lqb = JQA & ~JRB & ~KQA | ~JQA & JRB & ~KQA | ~JQA & ~JRB & KQA | ~JQA & ~JRB & ~KQA; 
	assign LRA = JRA & ~JSB & ~KRA | ~JRA & JSB & ~KRA | ~JRA & ~JSB & KRA | JRA & JSB & KRA; 
	assign lrb = JRA & ~JSB & ~KRA | ~JRA & JSB & ~KRA | ~JRA & ~JSB & KRA | ~JRA & ~JSB & ~KRA; 
	assign LSA = JSA & ~JTB & ~KSA | ~JSA & JTB & ~KSA | ~JSA & ~JTB & KSA | JSA & JTB & KSA; 
	assign lsb = JSA & ~JTB & ~KSA | ~JSA & JTB & ~KSA | ~JSA & ~JTB & KSA | ~JSA & ~JTB & ~KSA; 
	assign LTA = JTA & ~JUB & ~KTA | ~JTA & JUB & ~KTA | ~JTA & ~JUB & KTA | JTA & JUB & KTA; 
	assign ltb = JTA & ~JUB & ~KTA | ~JTA & JUB & ~KTA | ~JTA & ~JUB & KTA | ~JTA & ~JUB & ~KTA; 
	assign LUA = JUA & ~JVB & ~KUA | ~JUA & JVB & ~KUA | ~JUA & ~JVB & KUA | JUA & JVB & KUA; 
	assign lub = JUA & ~JVB & ~KUA | ~JUA & JVB & ~KUA | ~JUA & ~JVB & KUA | ~JUA & ~JVB & ~KUA; 
	assign LVA = JVA & ~JWB & ~KVA | ~JVA & JWB & ~KVA | ~JVA & ~JWB & KVA | JVA & JWB & KVA; 
	assign lvb = JVA & ~JWB & ~KVA | ~JVA & JWB & ~KVA | ~JVA & ~JWB & KVA | ~JVA & ~JWB & ~KVA; 
	assign NHC = ~nee & NAF | ~nef; 
	assign NHD = ~nee & NAF & NAG | ~nef & NAG | ~neg; 
	assign NHE = ~nee & NAF & NAG & NAH | ~nef & NAG & NAH | ~neg & NAH | NEH; 
	assign NIC = ~nei & NAJ | ~nej; 
	assign NID = ~nei & NAJ & NAK | ~nej & NAK | ~nek; 
	assign NIE = ~nei & NAJ & NAK & NAL | ~nej & NAK & NAL | ~nek & NAL | ~nel; 
	assign NJC = ~nem & NAN | ~nen; 
	assign NJD = ~nem & NAN & NAO | ~nen & NAO | ~neo; 
	assign NJE = ~nem & NAN & NAO & NAP | ~nen & NAO & NAP | ~neo & NAP | ~nep; 
	assign NKC = ~nfa & NBB | ~nfb; 
	assign NKD = ~nfa & NBB & NBC | ~nfb & NBC | ~nfc; 
	assign NKE = ~nfa & NBB & NBC & NBD | ~nfb & NBC & NBD | ~nfc & NBD | ~nfd; 
	assign NLC = ~nfe & NBF | ~nff; 
	assign NLD = ~nfe & NBF & NBG | ~nff & NBG | ~nfg; 
	assign NLE = ~nfe & NBF & NBG & NBH | ~nff & NBG & NBH | ~nfg & NBH | ~nfh; 
	assign ENC = ~dkh & ~DKJ | dkh & DKJ; 
	assign CIE = BAI & ACI; 
	assign CIF = BAI & ACK; 
	assign CIG = BAI & ACM; 
	assign CIH = BAI & ACO; 
	assign CII = BAI & ADA; 
	assign CIJ = BAI & ADC; 
	assign CIK = BAI & ADE; 
	assign CIL = BAI & ADG; 
	assign CJA = BAJ & ACQ; 
	assign CJB = BAJ & ACB; 
	assign CJC = BAJ & ACD; 
	assign CJD = BAJ & ACF; 
	assign CJE = BAJ & ACH; 
	assign CJF = BAJ & ACJ; 
	assign CJG = BAJ & ACL; 
	assign CJH = BAJ & ACN; 
	assign CJI = BAJ & ACP; 
	assign CJJ = BAJ & ADB; 
	assign CJK = BAJ & ADD; 
	assign CJL = BAJ & ADF; 
	assign CKA = BAK & ACA; 
	assign NMC = ~nfi & NBJ | ~nfj; 
	assign NMD = ~nfi & NBJ & NBK | ~nfj & NBK | ~nfk; 
	assign CKB = BAK & ACC; 
	assign CKC = BAK & ACE; 
	assign CKD = BAK & ACG; 
	assign NME = ~nfi & NBJ & NBK & NBL | ~nfj & NBK & NBL | ~nfk & NBL | ~nfl; 
	assign LWA = JWA & ~JXB & ~KWA | ~JWA & JXB & ~KWA | ~JWA & ~JXB & KWA | JWA & JXB & KWA; 
	assign lwb = JWA & ~JXB & ~KWA | ~JWA & JXB & ~KWA | ~JWA & ~JXB & KWA | ~JWA & ~JXB & ~KWA; 
	assign LXA = JXA & ~JYB & ~KXA | ~JXA & JYB & ~KXA | ~JXA & ~JYB & KXA | JXA & JYB & KXA; 
	assign lxb = JXA & ~JYB & ~KXA | ~JXA & JYB & ~KXA | ~JXA & ~JYB & KXA | ~JXA & ~JYB & ~KXA; 
	assign LYA = JYA & ~KYA | ~JYA & KYA; 
	assign LZA = JZA & ~KZA & ~JZD | ~JZA & KZA & ~JZD | ~JZA & ~KZA & JZD | JZA & KZA & JZD; 
	assign lzb = JZA & ~KZA & ~JZD | ~JZA & KZA & ~JZD | ~JZA & ~KZA & JZD | ~JZA & ~KZA & ~JZD; 
	assign LZF = JZE & ~KZE | ~JZE & KZE; 
	assign LZD = JZC & ~KZC & ~KZF | ~JZC & KZC & ~KZF | ~JZC & ~KZC & KZF | JZC & KZC & KZF; 
	assign lze = JZC & ~KZC & ~KZF | ~JZC & KZC & ~KZF | ~JZC & ~KZC & KZF | ~JZC & ~KZC & ~KZF; 
	assign LZH = JZG & ~KZG | ~JZG & KZG; 
	assign LZI = JZG & KZG; 
	assign LGD = KGA & ~khb; 
	assign NND = ~nfm & NBN & NBO | ~nfn & NBO | ~nfo; 
	assign NNE = ~nfm & NBN & NBO & NBP | ~nfn & NBO & NBP | ~nfo & NBP | ~nfp; 
	assign LZJ = JZI & ~KZI | ~JZI & KZI; 
	assign LZL = JZK & ~KZJ | ~JZK & KZJ; 
	assign NUD = NBI & NBJ & NBK | NBK & ~nfj | ~nfk; 
	assign LZM = JZK & KZJ; 
	assign LYB = JYA & KYA; 
	assign LZN = JZL & ~KZL | ~JZL & KZL; 
	assign LZO = JZL & KZL; 
	assign CKE = BAK & ACI; 
	assign CKF = BAK & ACK; 
	assign CKG = BAK & ACM; 
	assign HXA = GXA & ~GYB | ~GXA & GYB; 
	assign HXB = GXA & GYB; 
	assign HYB = GYA & GZB; 
	assign HYA = GYA & ~GZB | ~GYA & GZB; 
	assign CKH = BAK & ACO; 
	assign CKI = BAK & ADA; 
	assign CKJ = BAK & ADC; 
	assign CKK = BAK & ADE; 
	assign CLA = BAL & ACQ; 
	assign CLB = BAL & ACB; 
	assign LFD = KFC & ~kgb ; 
	assign LHC = ~KHC & ~kib ; 
	assign LIC = ~KHC & ~kjb ; 
	assign CLC = BAL & ACD; 
	assign CLD = BAL & ACF; 
	assign CLE = BAL & ACH; 
	assign CLF = BAL & ACJ; 
	assign CLG = BAL & ACL; 
	assign CLH = BAL & ACN; 
	assign CLI = BAL & ACP; 
	assign CLJ = BAL & ADB; 
	assign CLK = BAL & ADD; 
	assign CMA = BAM & ACA; 
	assign CMB = BAM & ACC; 
	assign CMC = BAM & ACE; 
	assign CMD = BAM & ACG; 
	assign CME = BAM & ACI; 
	assign CMF = BAM & ACK; 
	assign nxg = ~NBI | ~NBJ | ~NBK | ~NBL;
	assign nxi = ~NAE | ~NAF | ~NAG | ~NAH | ~NAI;
	assign nxj = ~NAJ | ~NAK | ~NAL | ~NAM | ~NAN;
	assign nxk = ~NAO | ~NAP | ~NBA | ~NBB | ~NBC;
	assign nxl = ~NBD | ~NBE | ~NBF | ~NBG | ~NBH;
	assign LHD = ~kib & KHC; 
	assign NUC = NBI & NBJ | ~nfj; 
	assign EUE = DOM & ~DOO | ~DOM & DOO; 
	assign CMG = BAM & ACM; 
	assign CMH = BAM & ACO; 
	assign CMI = BAM & ADA; 
	assign CMJ = BAM & ADC; 
	assign CNA = BAN & ACQ; 
	assign CNB = BAN & ACB; 
	assign LZG = JZE & KZE; 
	assign LZK = JZI & KZI; 
	assign CNC = BAN & ACD; 
	assign CND = BAN & ACF; 
	assign CNE = BAN & ACH; 
	assign NVC = NBM & NBN | ~nfn; 
	assign CNF = BAN & ACJ; 
	assign CNG = BAN & ACL; 
	assign CNH = BAN & ACN; 
	assign NVD = NBM & NBN & NBO | NBO & ~nfn | ~nfo; 
	assign CNI = BAN & ACP; 
	assign CNJ = BAN & ADB; 
	assign COA = BAO & ACA; 
	assign NRD = NAM & NAN & NAO | NAO & ~nen | ~neo; 
	assign NRC = NAM & NAN | ~nen; 
	assign COB = BAO & ACC; 
	assign COC = BAO & ACE; 
	assign COD = BAO & ACG; 
	assign COE = BAO & ACI; 
	assign COF = BAO & ACK; 
	assign COG = BAO & ACM; 
	assign FFH = DTS & DTU; 
	assign EMD = DKG & DKI; 
	assign EFB = ~dgh & ~dgk; 
	assign EEB = DGG & DGJ; 
	assign ECB = DGD & DGF; 
	assign COH = BAO & ACO; 
	assign COI = BAO & ADA; 
	assign CPA = BAP & ACQ; 
  	
	always@(posedge IZZ )
		begin 
			AAA <= IAA & ~QAA | AAB & QAA; 
			AAB <= IAB & ~QAA | AAC & QAA; 
			AAC <= IAC & ~QAA | AAD & QAA; 
			AAD <= IAD & ~QAA | AAE & QAA; 
			AAE <= IAE & ~QAA | AAF & QAA; 
			AAF <= IAF & ~QAA | AAG & QAA; 
			AAG <= IAG & ~QAA | AAH & QAA; 
			AAH <= IAH & ~QAA | AAI & QAA; 
			AAI <= IAI & ~QAA | AAJ & QAA; 
			AAJ <= IAJ & ~QAA | AAK & QAA; 
			AAK <= IAK & ~QAA | AAL & QAA; 
			AAL <= IAL & ~QAA | AAM & QAA; 
			AAM <= IAM & ~QAA | AAN & QAA; 
			AAN <= IAN & ~QAA | AAO & QAA; 
			AAO <= IAO & ~QAA | AAP & QAA; 
			AAP <= IAP & ~QAA | ABA & QAA; 
			AAQ <= QAA & AAA; 
			ABA <= IBA & ~QAA | ABB & QAA; 
			ABB <= IBB & ~QAA | ABC & QAA; 
			ABC <= IBC & ~QAA | ABD & QAA; 
			ABD <= IBD & ~QAA | ABE & QAA; 
			ABE <= IBE & ~QAA | ABF & QAA; 
			ABF <= IBF & ~QAA | ABG & QAA; 
			ABG <= IBG & ~QAA | ABH & QAA; 
			ABH <= IBH & ~QAA | ABI & QAA; 
			ABI <= IBI & ~QAA | ABJ & QAA; 
			ABJ <= IBJ & ~QAA | ABK & QAA; 
			ABK <= IBK & ~QAA | ABL & QAA; 
			ABL <= IBL & ~QAA | ABM & QAA; 
			ABM <= IBM & ~QAA | ABN & QAA; 
			ABN <= IBN & ~QAA | ABO & QAA; 
			ABO <= IBO & ~QAA | ABP & QAA; 
			ABP <= IBP & ~QAA | ZZO & QAA; 
			ACA <= AAA; 
			ACB <= AAB; 
			ACC <= AAC; 
			ACD <= AAD; 
			ACE <= AAE; 
			ACF <= AAF; 
			ACG <= AAG; 
			ACH <= AAH; 
			ACI <= AAI; 
			ACJ <= AAJ; 
			ACK <= AAK; 
			ACL <= AAL; 
			ACM <= AAM; 
			ACN <= AAN; 
			ACO <= AAO; 
			ACP <= AAP; 
			ACQ <= AAQ; 
			ADA <= ABA; 
			ADB <= ABB; 
			ADC <= ABC; 
			ADD <= ABD; 
			ADE <= ABE; 
			ADF <= ABF; 
			ADG <= ABG; 
			ADH <= ABH; 
			ADI <= ABI; 
			ADJ <= ABJ; 
			ADK <= ABK; 
			ADL <= ABL; 
			ADM <= ABM; 
			ADN <= ABN; 
			ADO <= ABO; 
			ADP <= ABP; 
			BAA <= IAA & ~QAB | BAA & QAB; 
			BAB <= IAB & ~QAB | BAB & QAB; 
			BAC <= IAC & ~QAB | BAC & QAB; 
			BAD <= IAD & ~QAB | BAD & QAB; 
			BAE <= IAE & ~QAB | BAE & QAB; 
			BAF <= IAF & ~QAB | BAF & QAB; 
			BAG <= IAG & ~QAB | BAG & QAB; 
			BAH <= IAH & ~QAB | BAH & QAB; 
			BAI <= IAI & ~QAB | BAI & QAB; 
			BAJ <= IAJ & ~QAB | BAJ & QAB; 
			BAK <= IAK & ~QAB | BAK & QAB; 
			BAL <= IAL & ~QAB | BAL & QAB; 
			BAM <= IAM & ~QAB | BAM & QAB; 
			BAN <= IAN & ~QAB | BAN & QAB; 
			BAO <= IAO & ~QAB | BAO & QAB; 
			BAP <= IAP & ~QAB | BAP & QAB; 
			BBA <= IBA & ~QAB | BBA & QAB; 
			BBB <= IBB & ~QAB | BBB & QAB; 
			BBC <= IBC & ~QAB | BBC & QAB; 
			BBD <= IBD & ~QAB | BBD & QAB; 
			BBE <= IBE & ~QAB | BBE & QAB; 
			BBF <= IBF & ~QAB | BBF & QAB; 
			BBG <= IBG & ~QAB | BBG & QAB; 
			BBH <= IBH & ~QAB | BBH & QAB; 
			BBI <= IBI & ~QAB | BBI & QAB; 
			BBJ <= IBJ & ~QAB | BBJ & QAB; 
			BBK <= IBK & ~QAB | BBK & QAB; 
			BBL <= ~QAB & IBL; 
			BBM <= ~QAB & IBM; 
			BBN <= ~QAB & IBN; 
			BBO <= IBO & ~QAB | BBO & QAB; 
			BBP <= IBP & ~QAB | BBP & QAB; 
			DGA <= CAA & ~CBA | ~CAA & CBA; 
			DGC <= CBA & CAA; 
			DGD <= CAB & ~CBB & ~CCA | ~CAB & CBB & ~CCA | ~CAB & ~CBB & CCA | CAB & CBB & CCA;
			dge <= CAB & ~CBB & ~CCA | ~CAB & CBB & ~CCA | ~CAB & ~CBB & CCA | ~CAB & ~CBB & ~CCA;
			DGF <= CDA; 
			DGG <= CAC & ~CBC & ~CCB | ~CAC & CBC & ~CCB | ~CAC & ~CBC & CCB | CAC & CBC & CCB;
			dgh <= CAC & ~CBC & ~CCB | ~CAC & CBC & ~CCB | ~CAC & ~CBC & CCB | ~CAC & ~CBC & ~CCB;
			DGJ <= CDB & ~CEA & ~CFA | ~CDB & CEA & ~CFA | ~CDB & ~CEA & CFA | CDB & CEA & CFA;
			dgk <= CDB & ~CEA & ~CFA | ~CDB & CEA & ~CFA | ~CDB & ~CEA & CFA | ~CDB & ~CEA & ~CFA;
			DHA <= CAD & ~CBD & ~CCC | ~CAD & CBD & ~CCC | ~CAD & ~CBD & CCC | CAD & CBD & CCC;
			dhb <= CAD & ~CBD & ~CCC | ~CAD & CBD & ~CCC | ~CAD & ~CBD & CCC | ~CAD & ~CBD & ~CCC;
			DHC <= CDC & ~CEB & ~CFB | ~CDC & CEB & ~CFB | ~CDC & ~CEB & CFB | CDC & CEB & CFB;
			dhd <= CDC & ~CEB & ~CFB | ~CDC & CEB & ~CFB | ~CDC & ~CEB & CFB | ~CDC & ~CEB & ~CFB;
			DHE <= CGA & ~CHA | ~CGA & CHA; 
			DHF <= CGA & CHA; 
			DIA <= CAE & ~CBE & ~CCD | ~CAE & CBE & ~CCD | ~CAE & ~CBE & CCD | CAE & CBE & CCD;
			dib <= CAE & ~CBE & ~CCD | ~CAE & CBE & ~CCD | ~CAE & ~CBE & CCD | ~CAE & ~CBE & ~CCD;
			DIC <= CDD & ~CEC & ~CFC | ~CDD & CEC & ~CFC | ~CDD & ~CEC & CFC | CDD & CEC & CFC;
			did <= CDD & ~CEC & ~CFC | ~CDD & CEC & ~CFC | ~CDD & ~CEC & CFC | ~CDD & ~CEC & ~CFC;
			DIE <= CGB & ~CHB & ~CIA | ~CGB & CHB & ~CIA | ~CGB & ~CHB & CIA | CGB & CHB & CIA;
			dif <= CGB & ~CHB & ~CIA | ~CGB & CHB & ~CIA | ~CGB & ~CHB & CIA | ~CGB & ~CHB & ~CIA;
			DIG <= CJA; 
			DJA <= CAF & ~CBF & ~CCE | ~CAF & CBF & ~CCE | ~CAF & ~CBF & CCE | CAF & CBF & CCE;
			djb <= CAF & ~CBF & ~CCE | ~CAF & CBF & ~CCE | ~CAF & ~CBF & CCE | ~CAF & ~CBF & ~CCE;
			DJC <= CDE & ~CED & ~CFD | ~CDE & CED & ~CFD | ~CDE & ~CED & CFD | CDE & CED & CFD;
			djd <= CDE & ~CED & ~CFD | ~CDE & CED & ~CFD | ~CDE & ~CED & CFD | ~CDE & ~CED & ~CFD;
			DJE <= CGC & ~CHC & ~CIB | ~CGC & CHC & ~CIB | ~CGC & ~CHC & CIB | CGC & CHC & CIB;
			djf <= CGC & ~CHC & ~CIB | ~CGC & CHC & ~CIB | ~CGC & ~CHC & CIB | ~CGC & ~CHC & ~CIB;
			DJG <= CJB & ~CKA & ~CLA | ~CJB & CKA & ~CLA | ~CJB & ~CKA & CLA | CJB & CKA & CLA;
			djh <= CJB & ~CKA & ~CLA | ~CJB & CKA & ~CLA | ~CJB & ~CKA & CLA | ~CJB & ~CKA & ~CLA;
			DKA <= CAG & ~CBG & ~CCF | ~CAG & CBG & ~CCF | ~CAG & ~CBG & CCF | CAG & CBG & CCF;
			dkb <= CAG & ~CBG & ~CCF | ~CAG & CBG & ~CCF | ~CAG & ~CBG & CCF | ~CAG & ~CBG & ~CCF;
			DKC <= CDF & ~CEE & ~CFE | ~CDF & CEE & ~CFE | ~CDF & ~CEE & CFE | CDF & CEE & CFE;
			dkd <= CDF & ~CEE & ~CFE | ~CDF & CEE & ~CFE | ~CDF & ~CEE & CFE | ~CDF & ~CEE & ~CFE;
			DKE <= CGD & ~CHD & ~CIC | ~CGD & CHD & ~CIC | ~CGD & ~CHD & CIC | CGD & CHD & CIC;
			dkf <= CGD & ~CHD & ~CIC | ~CGD & CHD & ~CIC | ~CGD & ~CHD & CIC | ~CGD & ~CHD & ~CIC;
			DKG <= CJC & ~CKB & ~CLB | ~CJC & CKB & ~CLB | ~CJC & ~CKB & CLB | CJC & CKB & CLB;
			dkh <= CJC & ~CKB & ~CLB | ~CJC & CKB & ~CLB | ~CJC & ~CKB & CLB | ~CJC & ~CKB & ~CLB;
			DKI <= CNA & ~CMA | ~CNA & CMA; 
			DKJ <= CMA & CNA; 
			DLA <= CAH & ~CBH & ~CCG | ~CAH & CBH & ~CCG | ~CAH & ~CBH & CCG | CAH & CBH & CCG;
			dlb <= CAH & ~CBH & ~CCG | ~CAH & CBH & ~CCG | ~CAH & ~CBH & CCG | ~CAH & ~CBH & ~CCG;
			DLC <= CDG & ~CEF & ~CFF | ~CDG & CEF & ~CFF | ~CDG & ~CEF & CFF | CDG & CEF & CFF;
			dld <= CDG & ~CEF & ~CFF | ~CDG & CEF & ~CFF | ~CDG & ~CEF & CFF | ~CDG & ~CEF & ~CFF;
			DLE <= CGE & ~CHE & ~CID | ~CGE & CHE & ~CID | ~CGE & ~CHE & CID | CGE & CHE & CID;
			dlf <= CGE & ~CHE & ~CID | ~CGE & CHE & ~CID | ~CGE & ~CHE & CID | ~CGE & ~CHE & ~CID;
			DLG <= CJD & ~CKC & ~CLC | ~CJD & CKC & ~CLC | ~CJD & ~CKC & CLC | CJD & CKC & CLC;
			dlh <= CJD & ~CKC & ~CLC | ~CJD & CKC & ~CLC | ~CJD & ~CKC & CLC | ~CJD & ~CKC & ~CLC;
			DLI <= CMB & ~CNB & ~COA | ~CMB & CNB & ~COA | ~CMB & ~CNB & COA | CMB & CNB & COA;
			dlj <= CMB & ~CNB & ~COA | ~CMB & CNB & ~COA | ~CMB & ~CNB & COA | ~CMB & ~CNB & ~COA;
			DLK <= CPA; 
			DMA <= CAI & ~CBI & ~CCH | ~CAI & CBI & ~CCH | ~CAI & ~CBI & CCH | CAI & CBI & CCH;
			dmb <= CAI & ~CBI & ~CCH | ~CAI & CBI & ~CCH | ~CAI & ~CBI & CCH | ~CAI & ~CBI & ~CCH;
			DMC <= CDH & ~CEG & ~CFG | ~CDH & CEG & ~CFG | ~CDH & ~CEG & CFG | CDH & CEG & CFG;
			dmd <= CDH & ~CEG & ~CFG | ~CDH & CEG & ~CFG | ~CDH & ~CEG & CFG | ~CDH & ~CEG & ~CFG;
			DME <= CGF & ~CHF & ~CIE | ~CGF & CHF & ~CIE | ~CGF & ~CHF & CIE | CGF & CHF & CIE;
			dmf <= CGF & ~CHF & ~CIE | ~CGF & CHF & ~CIE | ~CGF & ~CHF & CIE | ~CGF & ~CHF & ~CIE;
			DMG <= CJE & ~CKD & ~CLD | ~CJE & CKD & ~CLD | ~CJE & ~CKD & CLD | CJE & CKD & CLD;
			dmh <= CJE & ~CKD & ~CLD | ~CJE & CKD & ~CLD | ~CJE & ~CKD & CLD | ~CJE & ~CKD & ~CLD;
			DMI <= CMC & ~CNC & ~COB | ~CMC & CNC & ~COB | ~CMC & ~CNC & COB | CMC & CNC & COB;
			dmj <= CMC & ~CNC & ~COB | ~CMC & CNC & ~COB | ~CMC & ~CNC & COB | ~CMC & ~CNC & ~COB;
			DMK <= CPB & ~CQA & ~CRA | ~CPB & CQA & ~CRA | ~CPB & ~CQA & CRA | CPB & CQA & CRA;
			dml <= CPB & ~CQA & ~CRA | ~CPB & CQA & ~CRA | ~CPB & ~CQA & CRA | ~CPB & ~CQA & ~CRA;
			DNA <= CAJ & ~CBJ & ~CCI | ~CAJ & CBJ & ~CCI | ~CAJ & ~CBJ & CCI | CAJ & CBJ & CCI;
			dnb <= CAJ & ~CBJ & ~CCI | ~CAJ & CBJ & ~CCI | ~CAJ & ~CBJ & CCI | ~CAJ & ~CBJ & ~CCI;
			DNC <= CDI & ~CEH & ~CFH | ~CDI & CEH & ~CFH | ~CDI & ~CEH & CFH | CDI & CEH & CFH;
			dnd <= CDI & ~CEH & ~CFH | ~CDI & CEH & ~CFH | ~CDI & ~CEH & CFH | ~CDI & ~CEH & ~CFH;
			DNE <= CGG & ~CHG & ~CIF | ~CGG & CHG & ~CIF | ~CGG & ~CHG & CIF | CGG & CHG & CIF;
			dnf <= CGG & ~CHG & ~CIF | ~CGG & CHG & ~CIF | ~CGG & ~CHG & CIF | ~CGG & ~CHG & ~CIF;
			DNG <= CJF & ~CKE & ~CLE | ~CJF & CKE & ~CLE | ~CJF & ~CKE & CLE | CJF & CKE & CLE;
			dnh <= CJF & ~CKE & ~CLE | ~CJF & CKE & ~CLE | ~CJF & ~CKE & CLE | ~CJF & ~CKE & ~CLE;
			DNI <= CMD & ~CND & ~COC | ~CMD & CND & ~COC | ~CMD & ~CND & COC | CMD & CND & COC;
			dnj <= CMD & ~CND & ~COC | ~CMD & CND & ~COC | ~CMD & ~CND & COC | ~CMD & ~CND & ~COC;
			DNK <= CPC & ~CQB & ~CRB | ~CPC & CQB & ~CRB | ~CPC & ~CQB & CRB | CPC & CQB & CRB;
			dnl <= CPC & ~CQB & ~CRB | ~CPC & CQB & ~CRB | ~CPC & ~CQB & CRB | ~CPC & ~CQB & ~CRB;
			DNM <= CSA & ~CTA | ~CSA & CTA; 
			DNO <= CTA & CSA; 
			DOA <= CAK & ~CBK & ~CCJ | ~CAK & CBK & ~CCJ | ~CAK & ~CBK & CCJ | CAK & CBK & CCJ;
			dob <= CAK & ~CBK & ~CCJ | ~CAK & CBK & ~CCJ | ~CAK & ~CBK & CCJ | ~CAK & ~CBK & ~CCJ;
			DOC <= CDJ & ~CEI & ~CFI | ~CDJ & CEI & ~CFI | ~CDJ & ~CEI & CFI | CDJ & CEI & CFI;
			dod <= CDJ & ~CEI & ~CFI | ~CDJ & CEI & ~CFI | ~CDJ & ~CEI & CFI | ~CDJ & ~CEI & ~CFI;
			DOE <= CGH & ~CHH & ~CIG | ~CGH & CHH & ~CIG | ~CGH & ~CHH & CIG | CGH & CHH & CIG;
			dof <= CGH & ~CHH & ~CIG | ~CGH & CHH & ~CIG | ~CGH & ~CHH & CIG | ~CGH & ~CHH & ~CIG;
			DOG <= CJG & ~CKF & ~CLF | ~CJG & CKF & ~CLF | ~CJG & ~CKF & CLF | CJG & CKF & CLF;
			doh <= CJG & ~CKF & ~CLF | ~CJG & CKF & ~CLF | ~CJG & ~CKF & CLF | ~CJG & ~CKF & ~CLF;
			DOI <= CME & ~CNE & ~COD | ~CME & CNE & ~COD | ~CME & ~CNE & COD | CME & CNE & COD;
			doj <= CME & ~CNE & ~COD | ~CME & CNE & ~COD | ~CME & ~CNE & COD | ~CME & ~CNE & ~COD;
			DOK <= CPD & ~CQC & ~CRC | ~CPD & CQC & ~CRC | ~CPD & ~CQC & CRC | CPD & CQC & CRC;
			dol <= CPD & ~CQC & ~CRC | ~CPD & CQC & ~CRC | ~CPD & ~CQC & CRC | ~CPD & ~CQC & ~CRC;
			DOM <= CSB & ~CTB & ~CUA | ~CSB & CTB & ~CUA | ~CSB & ~CTB & CUA | CSB & CTB & CUA;
			don <= CSB & ~CTB & ~CUA | ~CSB & CTB & ~CUA | ~CSB & ~CTB & CUA | ~CSB & ~CTB & ~CUA;
			DOO <= CVA; 
			DPA <= CAL & ~CBL & ~CCK | ~CAL & CBL & ~CCK | ~CAL & ~CBL & CCK | CAL & CBL & CCK;
			dpb <= CAL & ~CBL & ~CCK | ~CAL & CBL & ~CCK | ~CAL & ~CBL & CCK | ~CAL & ~CBL & ~CCK;
			DPC <= CDK & ~CEJ & ~CFJ | ~CDK & CEJ & ~CFJ | ~CDK & ~CEJ & CFJ | CDK & CEJ & CFJ;
			dpd <= CDK & ~CEJ & ~CFJ | ~CDK & CEJ & ~CFJ | ~CDK & ~CEJ & CFJ | ~CDK & ~CEJ & ~CFJ;
			DPE <= CGI & ~CHI & ~CIH | ~CGI & CHI & ~CIH | ~CGI & ~CHI & CIH | CGI & CHI & CIH;
			dpf <= CGI & ~CHI & ~CIH | ~CGI & CHI & ~CIH | ~CGI & ~CHI & CIH | ~CGI & ~CHI & ~CIH;
			DPG <= CJH & ~CKG & ~CLG | ~CJH & CKG & ~CLG | ~CJH & ~CKG & CLG | CJH & CKG & CLG;
			dph <= CJH & ~CKG & ~CLG | ~CJH & CKG & ~CLG | ~CJH & ~CKG & CLG | ~CJH & ~CKG & ~CLG;
			DPI <= CMF & ~CNF & ~COE | ~CMF & CNF & ~COE | ~CMF & ~CNF & COE | CMF & CNF & COE;
			dpj <= CMF & ~CNF & ~COE | ~CMF & CNF & ~COE | ~CMF & ~CNF & COE | ~CMF & ~CNF & ~COE;
			DPK <= CPE & ~CQD & ~CRD | ~CPE & CQD & ~CRD | ~CPE & ~CQD & CRD | CPE & CQD & CRD;
			dpl <= CPE & ~CQD & ~CRD | ~CPE & CQD & ~CRD | ~CPE & ~CQD & CRD | ~CPE & ~CQD & ~CRD;
			DPM <= CSC & ~CTC & ~CUB | ~CSC & CTC & ~CUB | ~CSC & ~CTC & CUB | CSC & CTC & CUB;
			dpn <= CSC & ~CTC & ~CUB | ~CSC & CTC & ~CUB | ~CSC & ~CTC & CUB | ~CSC & ~CTC & ~CUB;
			DPO <= CVB & ~CWA & ~CXA | ~CVB & CWA & ~CXA | ~CVB & ~CWA & CXA | CVB & CWA & CXA;
			dpp <= CVB & ~CWA & ~CXA | ~CVB & CWA & ~CXA | ~CVB & ~CWA & CXA | ~CVB & ~CWA & ~CXA;
			DQA <= CAM & ~CBM & ~CCL | ~CAM & CBM & ~CCL | ~CAM & ~CBM & CCL | CAM & CBM & CCL;
			dqb <= CAM & ~CBM & ~CCL | ~CAM & CBM & ~CCL | ~CAM & ~CBM & CCL | ~CAM & ~CBM & ~CCL;
			DQC <= CDL & ~CEK & ~CFK | ~CDL & CEK & ~CFK | ~CDL & ~CEK & CFK | CDL & CEK & CFK;
			dqd <= CDL & ~CEK & ~CFK | ~CDL & CEK & ~CFK | ~CDL & ~CEK & CFK | ~CDL & ~CEK & ~CFK;
			DQE <= CGJ & ~CHJ & ~CII | ~CGJ & CHJ & ~CII | ~CGJ & ~CHJ & CII | CGJ & CHJ & CII;
			dqf <= CGJ & ~CHJ & ~CII | ~CGJ & CHJ & ~CII | ~CGJ & ~CHJ & CII | ~CGJ & ~CHJ & ~CII;
			DQG <= CJI & ~CKH & ~CLH | ~CJI & CKH & ~CLH | ~CJI & ~CKH & CLH | CJI & CKH & CLH;
			dqh <= CJI & ~CKH & ~CLH | ~CJI & CKH & ~CLH | ~CJI & ~CKH & CLH | ~CJI & ~CKH & ~CLH;
			DQI <= CMG & ~CNG & ~COF | ~CMG & CNG & ~COF | ~CMG & ~CNG & COF | CMG & CNG & COF;
			dqj <= CMG & ~CNG & ~COF | ~CMG & CNG & ~COF | ~CMG & ~CNG & COF | ~CMG & ~CNG & ~COF;
			DQK <= CPF & ~CQE & ~CRE | ~CPF & CQE & ~CRE | ~CPF & ~CQE & CRE | CPF & CQE & CRE;
			dql <= CPF & ~CQE & ~CRE | ~CPF & CQE & ~CRE | ~CPF & ~CQE & CRE | ~CPF & ~CQE & ~CRE;
			DQM <= CSD & ~CTD & ~CUC | ~CSD & CTD & ~CUC | ~CSD & ~CTD & CUC | CSD & CTD & CUC;
			dqn <= CSD & ~CTD & ~CUC | ~CSD & CTD & ~CUC | ~CSD & ~CTD & CUC | ~CSD & ~CTD & ~CUC;
			DQO <= CVC & ~CWB & ~CXB | ~CVC & CWB & ~CXB | ~CVC & ~CWB & CXB | CVC & CWB & CXB;
			dqp <= CVC & ~CWB & ~CXB | ~CVC & CWB & ~CXB | ~CVC & ~CWB & CXB | ~CVC & ~CWB & ~CXB;
			DQQ <= ~CZA & CYA; 
			DQR <= CZA & CYA; 
			DRA <= CAN & ~CBN & ~CCM | ~CAN & CBN & ~CCM | ~CAN & ~CBN & CCM | CAN & CBN & CCM;
			drb <= CAN & ~CBN & ~CCM | ~CAN & CBN & ~CCM | ~CAN & ~CBN & CCM | ~CAN & ~CBN & ~CCM;
			DRC <= CDM & ~CEL & ~CFL | ~CDM & CEL & ~CFL | ~CDM & ~CEL & CFL | CDM & CEL & CFL;
			drd <= CDM & ~CEL & ~CFL | ~CDM & CEL & ~CFL | ~CDM & ~CEL & CFL | ~CDM & ~CEL & ~CFL;
			DRE <= CGK & ~CHK & ~CIJ | ~CGK & CHK & ~CIJ | ~CGK & ~CHK & CIJ | CGK & CHK & CIJ;
			drf <= CGK & ~CHK & ~CIJ | ~CGK & CHK & ~CIJ | ~CGK & ~CHK & CIJ | ~CGK & ~CHK & ~CIJ;
			DRG <= CJJ & ~CKI & ~CLI | ~CJJ & CKI & ~CLI | ~CJJ & ~CKI & CLI | CJJ & CKI & CLI;
			drh <= CJJ & ~CKI & ~CLI | ~CJJ & CKI & ~CLI | ~CJJ & ~CKI & CLI | ~CJJ & ~CKI & ~CLI;
			DRI <= CMH & ~CNH & ~COG | ~CMH & CNH & ~COG | ~CMH & ~CNH & COG | CMH & CNH & COG;
			drj <= CMH & ~CNH & ~COG | ~CMH & CNH & ~COG | ~CMH & ~CNH & COG | ~CMH & ~CNH & ~COG;
			DRK <= CPG & ~CQF & ~CRF | ~CPG & CQF & ~CRF | ~CPG & ~CQF & CRF | CPG & CQF & CRF;
			drl <= CPG & ~CQF & ~CRF | ~CPG & CQF & ~CRF | ~CPG & ~CQF & CRF | ~CPG & ~CQF & ~CRF;
			DRM <= CSE & ~CTE & ~CUD | ~CSE & CTE & ~CUD | ~CSE & ~CTE & CUD | CSE & CTE & CUD;
			drn <= CSE & ~CTE & ~CUD | ~CSE & CTE & ~CUD | ~CSE & ~CTE & CUD | ~CSE & ~CTE & ~CUD;
			DRO <= CVD & ~CWC & ~CXC | ~CVD & CWC & ~CXC | ~CVD & ~CWC & CXC | CVD & CWC & CXC;
			drp <= CVD & ~CWC & ~CXC | ~CVD & CWC & ~CXC | ~CVD & ~CWC & CXC | ~CVD & ~CWC & ~CXC;
			DRQ <= CYB & ~CZB & ~DAA | ~CYB & CZB & ~DAA | ~CYB & ~CZB & DAA | CYB & CZB & DAA;
			drr <= CYB & ~CZB & ~DAA | ~CYB & CZB & ~DAA | ~CYB & ~CZB & DAA | ~CYB & ~CZB & ~DAA;
			DRS <= DBA; 
			DSA <= CAO & ~CBO & ~CCN | ~CAO & CBO & ~CCN | ~CAO & ~CBO & CCN | CAO & CBO & CCN;
			dsb <= CAO & ~CBO & ~CCN | ~CAO & CBO & ~CCN | ~CAO & ~CBO & CCN | ~CAO & ~CBO & ~CCN;
			DSC <= CDN & ~CEM & ~CFM | ~CDN & CEM & ~CFM | ~CDN & ~CEM & CFM | CDN & CEM & CFM;
			dsd <= CDN & ~CEM & ~CFM | ~CDN & CEM & ~CFM | ~CDN & ~CEM & CFM | ~CDN & ~CEM & ~CFM;
			DSE <= CGL & ~CHL & ~CIK | ~CGL & CHL & ~CIK | ~CGL & ~CHL & CIK | CGL & CHL & CIK;
			dsf <= CGL & ~CHL & ~CIK | ~CGL & CHL & ~CIK | ~CGL & ~CHL & CIK | ~CGL & ~CHL & ~CIK;
			DSG <= CJK & ~CKJ & ~CLJ | ~CJK & CKJ & ~CLJ | ~CJK & ~CKJ & CLJ | CJK & CKJ & CLJ;
			dsh <= CJK & ~CKJ & ~CLJ | ~CJK & CKJ & ~CLJ | ~CJK & ~CKJ & CLJ | ~CJK & ~CKJ & ~CLJ;
			DSI <= CMI & ~CNI & ~COH | ~CMI & CNI & ~COH | ~CMI & ~CNI & COH | CMI & CNI & COH;
			dsj <= CMI & ~CNI & ~COH | ~CMI & CNI & ~COH | ~CMI & ~CNI & COH | ~CMI & ~CNI & ~COH;
			DSK <= CPH & ~CQG & ~CRG | ~CPH & CQG & ~CRG | ~CPH & ~CQG & CRG | CPH & CQG & CRG;
			dsl <= CPH & ~CQG & ~CRG | ~CPH & CQG & ~CRG | ~CPH & ~CQG & CRG | ~CPH & ~CQG & ~CRG;
			DSM <= CSF & ~CTF & ~CUE | ~CSF & CTF & ~CUE | ~CSF & ~CTF & CUE | CSF & CTF & CUE;
			dsn <= CSF & ~CTF & ~CUE | ~CSF & CTF & ~CUE | ~CSF & ~CTF & CUE | ~CSF & ~CTF & ~CUE;
			DSO <= CVE & ~CWD & ~CXD | ~CVE & CWD & ~CXD | ~CVE & ~CWD & CXD | CVE & CWD & CXD;
			dsp <= CVE & ~CWD & ~CXD | ~CVE & CWD & ~CXD | ~CVE & ~CWD & CXD | ~CVE & ~CWD & ~CXD;
			DSQ <= CYC & ~CZC & ~DAB | ~CYC & CZC & ~DAB | ~CYC & ~CZC & DAB | CYC & CZC & DAB;
			dsr <= CYC & ~CZC & ~DAB | ~CYC & CZC & ~DAB | ~CYC & ~CZC & DAB | ~CYC & ~CZC & ~DAB;
			DSS <= DBB & ~DCA & ~DDA | ~DBB & DCA & ~DDA | ~DBB & ~DCA & DDA | DBB & DCA & DDA;
			dst <= DBB & ~DCA & ~DDA | ~DBB & DCA & ~DDA | ~DBB & ~DCA & DDA | ~DBB & ~DCA & ~DDA;
			DTA <= CAP & ~CBP & ~CCO | ~CAP & CBP & ~CCO | ~CAP & ~CBP & CCO | CAP & CBP & CCO;
			dtb <= CAP & ~CBP & ~CCO | ~CAP & CBP & ~CCO | ~CAP & ~CBP & CCO | ~CAP & ~CBP & ~CCO;
			DTC <= CDO & ~CEN & ~CFN | ~CDO & CEN & ~CFN | ~CDO & ~CEN & CFN | CDO & CEN & CFN;
			dtd <= CDO & ~CEN & ~CFN | ~CDO & CEN & ~CFN | ~CDO & ~CEN & CFN | ~CDO & ~CEN & ~CFN;
			DTE <= CGM & ~CHM & ~CIL | ~CGM & CHM & ~CIL | ~CGM & ~CHM & CIL | CGM & CHM & CIL;
			dtf <= CGM & ~CHM & ~CIL | ~CGM & CHM & ~CIL | ~CGM & ~CHM & CIL | ~CGM & ~CHM & ~CIL;
			DTG <= CJL & ~CKK & ~CLK | ~CJL & CKK & ~CLK | ~CJL & ~CKK & CLK | CJL & CKK & CLK;
			dth <= CJL & ~CKK & ~CLK | ~CJL & CKK & ~CLK | ~CJL & ~CKK & CLK | ~CJL & ~CKK & ~CLK;
			DTI <= CMJ & ~CNJ & ~COI | ~CMJ & CNJ & ~COI | ~CMJ & ~CNJ & COI | CMJ & CNJ & COI;
			dtj <= CMJ & ~CNJ & ~COI | ~CMJ & CNJ & ~COI | ~CMJ & ~CNJ & COI | ~CMJ & ~CNJ & ~COI;
			DTK <= CPI & ~CQH & ~CRH | ~CPI & CQH & ~CRH | ~CPI & ~CQH & CRH | CPI & CQH & CRH;
			dtl <= CPI & ~CQH & ~CRH | ~CPI & CQH & ~CRH | ~CPI & ~CQH & CRH | ~CPI & ~CQH & ~CRH;
			DTM <= CSG & ~CTG & ~CUF | ~CSG & CTG & ~CUF | ~CSG & ~CTG & CUF | CSG & CTG & CUF;
			dtn <= CSG & ~CTG & ~CUF | ~CSG & CTG & ~CUF | ~CSG & ~CTG & CUF | ~CSG & ~CTG & ~CUF;
			DTO <= CVF & ~CWE & ~CXE | ~CVF & CWE & ~CXE | ~CVF & ~CWE & CXE | CVF & CWE & CXE;
			dtp <= CVF & ~CWE & ~CXE | ~CVF & CWE & ~CXE | ~CVF & ~CWE & CXE | ~CVF & ~CWE & ~CXE;
			DTQ <= CYD & ~CZD & ~DAC | ~CYD & CZD & ~DAC | ~CYD & ~CZD & DAC | CYD & CZD & DAC;
			dtr <= CYD & ~CZD & ~DAC | ~CYD & CZD & ~DAC | ~CYD & ~CZD & DAC | ~CYD & ~CZD & ~DAC;
			DTS <= DBC & ~DCB & ~DDB | ~DBC & DCB & ~DDB | ~DBC & ~DCB & DDB | DBC & DCB & DDB;
			dtt <= DBC & ~DCB & ~DDB | ~DBC & DCB & ~DDB | ~DBC & ~DCB & DDB | ~DBC & ~DCB & ~DDB;
			DTU <= DEA & ~DFA | ~DEA & DFA; 
			DTV <= DFA & DEA; 
			GAA <= FGA & ~FGC & ~FGE | ~FGA & FGC & ~FGE | ~FGA & ~FGC & FGE | FGA & FGC & FGE;
			gab <= FGA & ~FGC & ~FGE | ~FGA & FGC & ~FGE | ~FGA & ~FGC & FGE | ~FGA & ~FGC & ~FGE;
			GAC <= FGG & ffb & ffd | ~FGG & ~ffb & ffd | ~FGG & ffb & ~ffd | FGG & ~ffb & ~ffd;
			gad <= FGG & ffb & ffd | ~FGG & ~ffb & ffd | ~FGG & ffb & ~ffd | ~FGG & ffb & ffd;
			GAE <= ~fff & ~FFH | fff & FFH; 
			GAF <= FFH & ~fff; 
			GBA <= FFA & ~FFC & ~FFE | ~FFA & FFC & ~FFE | ~FFA & ~FFC & FFE | FFA & FFC & FFE;
			gbb <= FFA & ~FFC & ~FFE | ~FFA & FFC & ~FFE | ~FFA & ~FFC & FFE | ~FFA & ~FFC & ~FFE;
			GBC <= FFG & feb & fed | ~FFG & ~feb & fed | ~FFG & feb & ~fed | FFG & ~feb & ~fed;
			gbd <= FFG & feb & fed | ~FFG & ~feb & fed | ~FFG & feb & ~fed | ~FFG & feb & fed;
			GBE <= ~fef; 
			GCA <= FEA & ~FEC & dst | ~FEA & FEC & dst | ~FEA & ~FEC & ~dst | FEA & FEC & ~dst;
			gcb <= FEA & ~FEC & dst | ~FEA & FEC & dst | ~FEA & ~FEC & ~dst | ~FEA & ~FEC & dst;
			GCC <= ~fdf & fdb & fdd | fdf & ~fdb & fdd | fdf & fdb & ~fdd | ~fdf & ~fdb & ~fdd;
			gcd <= ~fdf & fdb & fdd | fdf & ~fdb & fdd | fdf & fdb & ~fdd | fdf & fdb & fdd;
			GCE <= FEE; 
			GDA <= FDA & ~FDC & ~FDE | ~FDA & FDC & ~FDE | ~FDA & ~FDC & FDE | FDA & FDC & FDE;
			gdb <= FDA & ~FDC & ~FDE | ~FDA & FDC & ~FDE | ~FDA & ~FDC & FDE | ~FDA & ~FDC & ~FDE;
			GDC <= DSS & fcb & fcd | ~DSS & ~fcb & fcd | ~DSS & fcb & ~fcd | DSS & ~fcb & ~fcd;
			gdd <= DSS & fcb & fcd | ~DSS & ~fcb & fcd | ~DSS & fcb & ~fcd | ~DSS & fcb & fcd;
			GDE <= ~fcf; 
			GEA <= FCA & ~FCC & ~FCE | ~FCA & FCC & ~FCE | ~FCA & ~FCC & FCE | FCA & FCC & FCE;
			geb <= FCA & ~FCC & ~FCE | ~FCA & FCC & ~FCE | ~FCA & ~FCC & FCE | ~FCA & ~FCC & ~FCE;
			GEC <= ~fbb & fbd & fbf | fbb & ~fbd & fbf | fbb & fbd & ~fbf | ~fbb & ~fbd & ~fbf;
			ged <= ~fbb & fbd & fbf | fbb & ~fbd & fbf | fbb & fbd & ~fbf | fbb & fbd & fbf;
			GFA <= FBA & ~FBC & ~FBE | ~FBA & FBC & ~FBE | ~FBA & ~FBC & FBE | FBA & FBC & FBE;
			gfb <= FBA & ~FBC & ~FBE | ~FBA & FBC & ~FBE | ~FBA & ~FBC & FBE | ~FBA & ~FBC & ~FBE;
			GFC <= DRS & fab & fad | ~DRS & ~fab & fad | ~DRS & fab & ~fad | DRS & ~fab & ~fad;
			gfd <= DRS & fab & fad | ~DRS & ~fab & fad | ~DRS & fab & ~fad | ~DRS & fab & fad;
			GFE <= ~faf; 
			GGA <= FAA & ~FAC & ~FAE | ~FAA & FAC & ~FAE | ~FAA & ~FAC & FAE | FAA & FAC & FAE;
			ggb <= FAA & ~FAC & ~FAE | ~FAA & FAC & ~FAE | ~FAA & ~FAC & FAE | ~FAA & ~FAC & ~FAE;
			GGC <= ~eyb & eyd & eyf | eyb & ~eyd & eyf | eyb & eyd & ~eyf | ~eyb & ~eyd & ~eyf;
			ggd <= ~eyb & eyd & eyf | eyb & ~eyd & eyf | eyb & eyd & ~eyf | eyb & eyd & eyf;
			GHA <= EYA & ~EYC & ~EYE | ~EYA & EYC & ~EYE | ~EYA & ~EYC & EYE | EYA & EYC & EYE;
			ghb <= EYA & ~EYC & ~EYE | ~EYA & EYC & ~EYE | ~EYA & ~EYC & EYE | ~EYA & ~EYC & ~EYE;
			GHC <= DQR & exb & exd | ~DQR & ~exb & exd | ~DQR & exb & ~exd | DQR & ~exb & ~exd;
			ghd <= DQR & exb & exd | ~DQR & ~exb & exd | ~DQR & exb & ~exd | ~DQR & exb & exd;
			GHE <= EXF; 
			GIA <= EXA & ~EXC & ~EXE | ~EXA & EXC & ~EXE | ~EXA & ~EXC & EXE | EXA & EXC & EXE;
			gib <= EXA & ~EXC & ~EXE | ~EXA & EXC & ~EXE | ~EXA & ~EXC & EXE | ~EXA & ~EXC & ~EXE;
			GIC <= ~ewb & ewd & ~EWF | ewb & ~ewd & ~EWF | ewb & ewd & EWF | ~ewb & ~ewd & EWF;
			gid <= ~ewb & ewd & ~EWF | ewb & ~ewd & ~EWF | ewb & ewd & EWF | ewb & ewd & ~EWF;
			GJA <= EWA & ~EWC & ~EWE | ~EWA & EWC & ~EWE | ~EWA & ~EWC & EWE | EWA & EWC & EWE;
			gjb <= EWA & ~EWC & ~EWE | ~EWA & EWC & ~EWE | ~EWA & ~EWC & EWE | ~EWA & ~EWC & ~EWE;
			GJC <= ~evb & evd | evb & ~evd; 
			GJD <= ~evd & ~evb; 
			GKA <= EVA & ~EVC & don | ~EVA & EVC & don | ~EVA & ~EVC & ~don | EVA & EVC & ~don;
			gkb <= EVA & ~EVC & don | ~EVA & EVC & don | ~EVA & ~EVC & ~don | ~EVA & ~EVC & don;
			GKC <= ~eub & eud & ~EUF | eub & ~eud & ~EUF | eub & eud & EUF | ~eub & ~eud & EUF;
			gkd <= ~eub & eud & ~EUF | eub & ~eud & ~EUF | eub & eud & EUF | eub & eud & ~EUF;
			GLA <= EUA & ~EUC & ~EUE | ~EUA & EUC & ~EUE | ~EUA & ~EUC & EUE | EUA & EUC & EUE;
			glb <= EUA & ~EUC & ~EUE | ~EUA & EUC & ~EUE | ~EUA & ~EUC & EUE | ~EUA & ~EUC & ~EUE;
			GLC <= ~etb & etd | etb & ~etd; 
			GLD <= ~etd & ~etb; 
			GMA <= ETA & ~ETC & ~DNO | ~ETA & ETC & ~DNO | ~ETA & ~ETC & DNO | ETA & ETC & DNO;
			gmb <= ETA & ~ETC & ~DNO | ~ETA & ETC & ~DNO | ~ETA & ~ETC & DNO | ~ETA & ~ETC & ~DNO;
			GMC <= ~esb & esd | esb & ~esd; 
			GMD <= ~esd & ~esb; 
			GNA <= ESA & ~ESC & ~DNM | ~ESA & ESC & ~DNM | ~ESA & ~ESC & DNM | ESA & ESC & DNM;
			gnb <= ESA & ~ESC & ~DNM | ~ESA & ESC & ~DNM | ~ESA & ~ESC & DNM | ~ESA & ~ESC & ~DNM;
			GNC <= ~erb & erd | erb & ~erd; 
			GND <= ~erd & ~erb; 
			GOA <= ERA & ~ERC & eqb | ~ERA & ERC & eqb | ~ERA & ~ERC & ~eqb | ERA & ERC & ~eqb;
			gob <= ERA & ~ERC & eqb | ~ERA & ERC & eqb | ~ERA & ~ERC & ~eqb | ~ERA & ~ERC & eqb;
			GOC <= ~eqd; 
			GPA <= EQA & ~EQC & epb | ~EQA & EQC & epb | ~EQA & ~EQC & ~epb | EQA & EQC & ~epb;
			gpb <= EQA & ~EQC & epb | ~EQA & EQC & epb | ~EQA & ~EQC & ~epb | ~EQA & ~EQC & epb;
			GPC <= EPD; 
			GQA <= EPA & ~EPC & eob | ~EPA & EPC & eob | ~EPA & ~EPC & ~eob | EPA & EPC & ~eob;
			gqb <= EPA & ~EPC & eob | ~EPA & EPC & eob | ~EPA & ~EPC & ~eob | ~EPA & ~EPC & eob;
			GQC <= ~eod; 
			GRA <= EOA & ~EOC & enb | ~EOA & EOC & enb | ~EOA & ~EOC & ~enb | EOA & EOC & ~enb;
			grb <= EOA & ~EOC & enb | ~EOA & EOC & enb | ~EOA & ~EOC & ~enb | ~EOA & ~EOC & enb;
			GRC <= END; 
			GSA <= ENA & ~ENC & emb | ~ENA & ENC & emb | ~ENA & ~ENC & ~emb | ENA & ENC & ~emb;
			gsb <= ENA & ~ENC & emb | ~ENA & ENC & emb | ~ENA & ~ENC & ~emb | ~ENA & ~ENC & emb;
			GSC <= EMD; 
			GTA <= EMA & ~EMC & elb | ~EMA & EMC & elb | ~EMA & ~EMC & ~elb | EMA & EMC & ~elb;
			gtb <= EMA & ~EMC & elb | ~EMA & EMC & elb | ~EMA & ~EMC & ~elb | ~EMA & ~EMC & elb;
			GUA <= ELA & djh & ekb | ~ELA & ~djh & ekb | ~ELA & djh & ~ekb | ELA & ~djh & ~ekb;
			gub <= ELA & djh & ekb | ~ELA & ~djh & ekb | ~ELA & djh & ~ekb | ~ELA & djh & ekb;
			GVA <= EKA & ~DJG & ejb | ~EKA & DJG & ejb | ~EKA & ~DJG & ~ejb | EKA & DJG & ~ejb;
			gvb <= EKA & ~DJG & ejb | ~EKA & DJG & ejb | ~EKA & ~DJG & ~ejb | ~EKA & ~DJG & ejb;
			GWA <= EJA & eib | ~EJA & ~eib; 
			GWB <= ~eib & EJA; 
			GXA <= EIA & ~DIG & ehb | ~EIA & DIG & ehb | ~EIA & ~DIG & ~ehb | EIA & DIG & ~ehb;
			gxb <= EIA & ~DIG & ehb | ~EIA & DIG & ehb | ~EIA & ~DIG & ~ehb | ~EIA & ~DIG & ehb;
			GYA <= EHA & egb | ~EHA & ~egb; 
			GYB <= ~egb & EHA; 
			GZA <= EGA & ~EFB | ~EGA & EFB; 
			GZB <= EFB & EGA; 
			GZD <= EFA & ~EEB | ~EFA & EEB; 
			GZE <= EEB & EFA; 
			GZF <= EEA; 
			GZH <= ECA; 
			GZK <= DGC; 
			GZL <= DGA; 
			GZM <= ~dge & ~ECB | dge & ECB; 
			GZN <= ECB & ~dge; 
			JAA <= HAA & ~HAC & hbb | ~HAA & HAC & hbb | ~HAA & ~HAC & ~hbb | HAA & HAC & ~hbb;
			jab <= HAA & ~HAC & hbb | ~HAA & HAC & hbb | ~HAA & ~HAC & ~hbb | ~HAA & ~HAC & hbb;
			JAC <= HBD; 
			JBA <= HBA & ~HBC & hcb | ~HBA & HBC & hcb | ~HBA & ~HBC & ~hcb | HBA & HBC & ~hcb;
			jbb <= HBA & ~HBC & hcb | ~HBA & HBC & hcb | ~HBA & ~HBC & ~hcb | ~HBA & ~HBC & hcb;
			JBC <= HCE; 
			JCA <= HCA & ~HCD & hdb | ~HCA & HCD & hdb | ~HCA & ~HCD & ~hdb | HCA & HCD & ~hdb;
			jcb <= HCA & ~HCD & hdb | ~HCA & HCD & hdb | ~HCA & ~HCD & ~hdb | ~HCA & ~HCD & hdb;
			JCC <= HDD; 
			JDA <= HDA & ~HDC & heb | ~HDA & HDC & heb | ~HDA & ~HDC & ~heb | HDA & HDC & ~heb;
			jdb <= HDA & ~HDC & heb | ~HDA & HDC & heb | ~HDA & ~HDC & ~heb | ~HDA & ~HDC & heb;
			JEA <= HEA & gfd & hfb | ~HEA & ~gfd & hfb | ~HEA & gfd & ~hfb | HEA & ~gfd & ~hfb;
			jeb <= HEA & gfd & hfb | ~HEA & ~gfd & hfb | ~HEA & gfd & ~hfb | ~HEA & gfd & hfb;
			JEC <= HFD; 
			JFA <= HFA & ~HFC & hgb | ~HFA & HFC & hgb | ~HFA & ~HFC & ~hgb | HFA & HFC & ~hgb;
			jfb <= HFA & ~HFC & hgb | ~HFA & HFC & hgb | ~HFA & ~HFC & ~hgb | ~HFA & ~HFC & hgb;
			JGA <= HGA & ghd & hhb | ~HGA & ~ghd & hhb | ~HGA & ghd & ~hhb | HGA & ~ghd & ~hhb;
			jgb <= HGA & ghd & hhb | ~HGA & ~ghd & hhb | ~HGA & ghd & ~hhb | ~HGA & ghd & hhb;
			JGC <= HHD; 
			JHA <= HHA & ~HHC & hib | ~HHA & HHC & hib | ~HHA & ~HHC & ~hib | HHA & HHC & ~hib;
			jhb <= HHA & ~HHC & hib | ~HHA & HHC & hib | ~HHA & ~HHC & ~hib | ~HHA & ~HHC & hib;
			JIA <= HIA & ~GJD & hjb | ~HIA & GJD & hjb | ~HIA & ~GJD & ~hjb | HIA & GJD & ~hjb;
			jib <= HIA & ~GJD & hjb | ~HIA & GJD & hjb | ~HIA & ~GJD & ~hjb | ~HIA & ~GJD & hjb;
			JJA <= HJA & gkd & hkb | ~HJA & ~gkd & hkb | ~HJA & gkd & ~hkb | HJA & ~gkd & ~hkb;
			jjb <= HJA & gkd & hkb | ~HJA & ~gkd & hkb | ~HJA & gkd & ~hkb | ~HJA & gkd & hkb;
			JKA <= HKA & ~GLD & hlb | ~HKA & GLD & hlb | ~HKA & ~GLD & ~hlb | HKA & GLD & ~hlb;
			jkb <= HKA & ~GLD & hlb | ~HKA & GLD & hlb | ~HKA & ~GLD & ~hlb | ~HKA & ~GLD & hlb;
			JLA <= HLA & ~GMD & hmb | ~HLA & GMD & hmb | ~HLA & ~GMD & ~hmb | HLA & GMD & ~hmb;
			jlb <= HLA & ~GMD & hmb | ~HLA & GMD & hmb | ~HLA & ~GMD & ~hmb | ~HLA & ~GMD & hmb;
			JMA <= HMA & ~GND & hnb | ~HMA & GND & hnb | ~HMA & ~GND & ~hnb | HMA & GND & ~hnb;
			jmb <= HMA & ~GND & hnb | ~HMA & GND & hnb | ~HMA & ~GND & ~hnb | ~HMA & ~GND & hnb;
			JNA <= HNA & hob | ~HNA & ~hob; 
			JNB <= ~hob & HNA; 
			JOA <= HOA & hpb | ~HOA & ~hpb; 
			JOB <= ~hpb & HOA; 
			JPA <= HPA & hqb | ~HPA & ~hqb; 
			JPB <= ~hqb & HPA; 
			JQA <= HQA & hrb | ~HQA & ~hrb; 
			JQB <= ~hrb & HQA; 
			JRA <= HRA & hsb | ~HRA & ~hsb; 
			JRB <= ~hsb & HRA; 
			JSA <= HSA & ~HTB | ~HSA & HTB; 
			JSB <= HTB & HSA; 
			JTA <= HTA & ~HUB | ~HTA & HUB; 
			JTB <= HUB & HTA; 
			JUA <= HUA & ~HVB | ~HUA & HVB; 
			JUB <= HVB & HUA; 
			JVA <= HVA & ~HWB | ~HVA & HWB; 
			JVB <= HWB & HVA; 
			JWA <= HWA & ~HXB | ~HWA & HXB; 
			JWB <= HXB & HWA; 
			JXA <= HXA & ~HYB | ~HXA & HYB; 
			JXB <= HYB & HXA; 
			JYA <= HYA & ~HZB | ~HYA & HZB; 
			JYB <= HZB & HYA; 
			JZA <= HZA; 
			JZC <= GZD & ~HZF | ~GZD & HZF; 
			JZD <= HZF & GZD; 
			JZE <= HZE; 
			JZG <= GZM; 
			JZI <= GZH; 
			JZK <= GZK; 
			JZL <= GZL; 
			KBA <= JAA; 
			kbb <= jab; 
			KBC <= JAC; 
			KCA <= JBA; 
			kcb <= jbb; 
			KCC <= JBC; 
			KDA <= JCA; 
			kdb <= jcb; 
			KDC <= JCC; 
			KEA <= JDA; 
			keb <= jdb; *************************************************
			KFA <= JEA; 
			kfb <= jeb; 
			KFC <= JEC; 
			KGA <= JFA; 
			kgb <= jfb; 
			KHA <= JGA; 
			khb <= jgb; 
			KHC <= JGC; 
			KIA <= JHA; 
			kib <= jhb; 
			KJA <= JIA; 
			kjb <= jib; 
			KKA <= JJA; 
			kkb <= jjb; 
			KLA <= JKA; 
			klb <= jkb; 
			KMA <= JLA; 
			kmb <= jlb; 
			KNA <= JMA; 
			knb <= jmb; 
			KOA <= JNA; 
			KOB <= JNB; 
			KPA <= JOA; 
			KPB <= JOB; 
			KQA <= JPA; 
			KQB <= JPB; 
			KRA <= JQA; 
			KRB <= JQB; 
			KSA <= JRA; 
			KSB <= JRB; 
			KTA <= JSA; 
			KTB <= JSB; 
			KUA <= JTA; 
			KUB <= JTB; 
			KVA <= JUA; 
			KVB <= JUB; 
			KWA <= JVA; 
			KWB <= JVB; 
			KXA <= JWA; 
			KXB <= JWB; 
			KYA <= JXA; 
			KYB <= JXB; 
			KZA <= JYA; 
			KZB <= JYB; 
			KZC <= JZA; 
			KZE <= JZC; 
			KZF <= JZD; 
			KZG <= JZE; 
			KZI <= JZG; 
			KZJ <= JZI; 
			KZL <= JZK; 
			KZM <= JZL; 
			MAA <= LBA & ~LBC & lcb | ~LBA & LBC & lcb | ~LBA & ~LBC & ~lcb | LBA & LBC & ~lcb;
			MAB <= LCA & ~LCC & kdb | ~LCA & LCC & kdb | ~LCA & ~LCC & ~kdb | LCA & LCC & ~kdb;
			MAC <= LDA & ~LDC & leb | ~LDA & LDC & leb | ~LDA & ~LDC & ~leb | LDA & LDC & ~leb;
			MAD <= LEA & ~LEC & lfb | ~LEA & LEC & lfb | ~LEA & ~LEC & ~lfb | LEA & LEC & ~lfb;
			MAE <= LFA & ~LFC & lgb | ~LFA & LFC & lgb | ~LFA & ~LFC & ~lgb | LFA & LFC & ~lgb;
			MAF <= LGA & ~LGC & lhb | ~LGA & LGC & lhb | ~LGA & ~LGC & ~lhb | LGA & LGC & ~lhb;
			MAG <= LHA & ~LHC & lib | ~LHA & LHC & lib | ~LHA & ~LHC & ~lib | LHA & LHC & ~lib;
			MAH <= LIA & ~LIC & ljb | ~LIA & LIC & ljb | ~LIA & ~LIC & ~ljb | LIA & LIC & ~ljb;
			MAI <= LJA & kkb & lkb | ~LJA & ~kkb & lkb | ~LJA & kkb & ~lkb | LJA & ~kkb & ~lkb;
			MAJ <= LKA & klb & llb | ~LKA & ~klb & llb | ~LKA & klb & ~llb | LKA & ~klb & ~llb;
			MAK <= LLA & kmb & lmb | ~LLA & ~kmb & lmb | ~LLA & kmb & ~lmb | LLA & ~kmb & ~lmb;
			MAL <= LMA & knb & lnb | ~LMA & ~knb & lnb | ~LMA & knb & ~lnb | LMA & ~knb & ~lnb;
			MAM <= LNA & ~KOB & lob | ~LNA & KOB & lob | ~LNA & ~KOB & ~lob | LNA & KOB & ~lob;
			MAN <= LOA & ~KPB & lpb | ~LOA & KPB & lpb | ~LOA & ~KPB & ~lpb | LOA & KPB & ~lpb;
			MAO <= LPA & ~KQB & lqb | ~LPA & KQB & lqb | ~LPA & ~KQB & ~lqb | LPA & KQB & ~lqb;
			MAP <= LQA & ~KRB & lrb | ~LQA & KRB & lrb | ~LQA & ~KRB & ~lrb | LQA & KRB & ~lrb;
			MBA <= LRA & ~KSB & lsb | ~LRA & KSB & lsb | ~LRA & ~KSB & ~lsb | LRA & KSB & ~lsb;
			MBB <= LSA & ~KTB & ltb | ~LSA & KTB & ltb | ~LSA & ~KTB & ~ltb | LSA & KTB & ~ltb;
			MBC <= LTA & ~KUB & lub | ~LTA & KUB & lub | ~LTA & ~KUB & ~lub | LTA & KUB & ~lub;
			MBD <= LUA & ~KVB & lvb | ~LUA & KVB & lvb | ~LUA & ~KVB & ~lvb | LUA & KVB & ~lvb;
			MBE <= LVA & ~KWB & lwb | ~LVA & KWB & lwb | ~LVA & ~KWB & ~lwb | LVA & KWB & ~lwb;
			MBF <= LWA & ~KXB & lxb | ~LWA & KXB & lxb | ~LWA & ~KXB & ~lxb | LWA & KXB & ~lxb;
			MBG <= LXA & ~KYB & ~LYB | ~LXA & KYB & ~LYB | ~LXA & ~KYB & LYB | LXA & KYB & LYB;
			MBH <= LYA & ~KZB & lzb | ~LYA & KZB & lzb | ~LYA & ~KZB & ~lzb | LYA & KZB & ~lzb;
			MBI <= LZA & ~ZZO & lze | ~LZA & ZZO & lze | ~LZA & ~ZZO & ~lze | LZA & ZZO & ~lze;
			MBJ <= LZD; 
			MBK <= LZF; 
			MBL <= LZH; 
			MBM <= LZJ; 
			MBN <= LZL; 
			MBO <= LZN; 
			MBP <= KZM; 
			mcb <= LCA & ~LCC & kdb | ~LCA & LCC & kdb | ~LCA & ~LCC & ~kdb | ~LCA & ~LCC & kdb;
			mcc <= LDA & ~LDC & leb | ~LDA & LDC & leb | ~LDA & ~LDC & ~leb | ~LDA & ~LDC & leb;
			mcd <= LEA & ~LEC & lfb | ~LEA & LEC & lfb | ~LEA & ~LEC & ~lfb | ~LEA & ~LEC & lfb;
			mce <= LFA & ~LFC & lgb | ~LFA & LFC & lgb | ~LFA & ~LFC & ~lgb | ~LFA & ~LFC & lgb;
			mcf <= LGA & ~LGC & lhb | ~LGA & LGC & lhb | ~LGA & ~LGC & ~lhb | ~LGA & ~LGC & lhb;
			mcg <= LHA & ~LHC & lib | ~LHA & LHC & lib | ~LHA & ~LHC & ~lib | ~LHA & ~LHC & lib;
			mch <= LIA & ~LIC & ljb | ~LIA & LIC & ljb | ~LIA & ~LIC & ~ljb | ~LIA & ~LIC & ljb;
			mci <= LJA & kkb & lkb | ~LJA & ~kkb & lkb | ~LJA & kkb & ~lkb | ~LJA & kkb & lkb;
			mcj <= LKA & klb & llb | ~LKA & ~klb & llb | ~LKA & klb & ~llb | ~LKA & klb & llb;
			mck <= LLA & kmb & lmb | ~LLA & ~kmb & lmb | ~LLA & kmb & ~lmb | ~LLA & kmb & lmb;
			mcl <= LMA & knb & lnb | ~LMA & ~knb & lnb | ~LMA & knb & ~lnb | ~LMA & knb & lnb;
			mcm <= LNA & ~KOB & lob | ~LNA & KOB & lob | ~LNA & ~KOB & ~lob | ~LNA & ~KOB & lob;
			mcn <= LOA & ~KPB & lpb | ~LOA & KPB & lpb | ~LOA & ~KPB & ~lpb | ~LOA & ~KPB & lpb;
			mco <= LPA & ~KQB & lqb | ~LPA & KQB & lqb | ~LPA & ~KQB & ~lqb | ~LPA & ~KQB & lqb;
			mcp <= LQA & ~KRB & lrb | ~LQA & KRB & lrb | ~LQA & ~KRB & ~lrb | ~LQA & ~KRB & lrb;
			mda <= LRA & ~KSB & lsb | ~LRA & KSB & lsb | ~LRA & ~KSB & ~lsb | ~LRA & ~KSB & lsb;
			mdb <= LSA & ~KTB & ltb | ~LSA & KTB & ltb | ~LSA & ~KTB & ~ltb | ~LSA & ~KTB & ltb;
			mdc <= LTA & ~KUB & lub | ~LTA & KUB & lub | ~LTA & ~KUB & ~lub | ~LTA & ~KUB & lub;
			mdd <= LUA & ~KVB & lvb | ~LUA & KVB & lvb | ~LUA & ~KVB & ~lvb | ~LUA & ~KVB & lvb;
			mde <= LVA & ~KWB & lwb | ~LVA & KWB & lwb | ~LVA & ~KWB & ~lwb | ~LVA & ~KWB & lwb;
			mdf <= LWA & ~KXB & lxb | ~LWA & KXB & lxb | ~LWA & ~KXB & ~lxb | ~LWA & ~KXB & lxb;
			mdg <= LXA & ~KYB & ~LYB | ~LXA & KYB & ~LYB | ~LXA & ~KYB & LYB | ~LXA & ~KYB & ~LYB;
			mdh <= LYA & ~KZB & lzb | ~LYA & KZB & lzb | ~LYA & ~KZB & ~lzb | ~LYA & ~KZB & lzb;
			mdi <= LZA & ~ZZO & lze | ~LZA & ZZO & lze | ~LZA & ~ZZO & ~lze | ~LZA & ~ZZO & lze;
			MDJ <= LZG; 
			MDK <= LZI; 
			MDL <= LZK; 
			MDM <= LZM; 
			MEA <= ~lcd; 
			MEB <= LDB & ldd | ~LDB & ~ldd; 
			MEC <= LDB & ~ldd | ZZO & ldd; 
			MED <= LED; 
			MEE <= LGD; 
			MEF <= LFD; 
			MEH <= LHD; 
			NAA <= MBP; 
			NAB <= MBO; 
			NAC <= MBN; 
			NAD <= MBM & ~MDM | ~MBM & MDM; 
			NAE <= MBL & ~MDL | ~MBL & MDL; 
			NAF <= MBK & ~MDK | ~MBK & MDK; 
			NAG <= MBJ & ~MDJ | ~MBJ & MDJ; 
			NAH <= MBI; 
			NAI <= MBH; 
			NAJ <= MBG & mdh | ~MBG & ~mdh; 
			NAK <= MBF & mdg | ~MBF & ~mdg; 
			NAL <= MBE & mdf | ~MBE & ~mdf; 
			NAM <= MBD & mde | ~MBD & ~mde; 
			NAN <= MBC & mdd | ~MBC & ~mdd; 
			NAO <= MBB & mdc | ~MBB & ~mdc; 
			NAP <= MBA & mdb | ~MBA & ~mdb; 
			NBA <= MAP & mda | ~MAP & ~mda; 
			NBB <= MAO & mcp | ~MAO & ~mcp; 
			NBC <= MAN & mco | ~MAN & ~mco; 
			NBD <= MAM & mcn | ~MAM & ~mcn; 
			NBE <= MAL & mcm | ~MAL & ~mcm; 
			NBF <= MAK & mcl | ~MAK & ~mcl; 
			NBG <= MAJ & mck | ~MAJ & ~mck; 
			NBH <= MAI & mcj | ~MAI & ~mcj; 
			NBI <= MAH & mci | ~MAH & ~mci; 
			NBJ <= MAG & mch | ~MAG & ~mch; 
			NBK <= MAF & mcg & ~MEH | ~MAF & ~mcg & ~MEH | ~MAF & mcg & MEH | MAF & ~mcg & MEH;
			NBL <= MAE & mcf & ~MEE | ~MAE & ~mcf & ~MEE | ~MAE & mcf & MEE | MAE & ~mcf & MEE;
			NBM <= MAD & mce & ~MEF | ~MAD & ~mce & ~MEF | ~MAD & mce & MEF | MAD & ~mce & MEF;
			NBN <= MAC & mcd & ~MED | ~MAC & ~mcd & ~MED | ~MAC & mcd & MED | MAC & ~mcd & MED;
			NBO <= MAB & mcc & ~MEB | ~MAB & ~mcc & ~MEB | ~MAB & mcc & MEB | MAB & ~mcc & MEB;
			NBP <= MAA & mcb & ~MEA | ~MAA & ~mcb & ~MEA | ~MAA & mcb & MEA | MAA & ~mcb & MEA;
			NED <= MBM & MDM; 
			nee <= ~MBL | ~MDL; 
			nef <= ~MBK | ~MDK; 
			neg <= ~MBJ | ~MDJ; 
			NEH <= ~mdi; 
			nei <= ~MBH | mdi; 
			nej <= ~MBG | mdh; 
			nek <= ~MBF | mdg; 
			nel <= ~MBE | mdf; 
			nem <= ~MBD | mde; 
			nen <= ~MBC | mdd; 
			neo <= ~MBB | mdc; 
			nep <= ~MBA | mdb; 
			nfa <= ~MAP | mda; 
			nfb <= ~MAO | mcp; 
			nfc <= ~MAN | mco; 
			nfd <= ~MAM | mcn; 
			nfe <= ~MAL | mcm; 
			nff <= ~MAK | mcl; 
			nfg <= ~MAJ | mck; 
			nfh <= ~MAI | mcj; 
			nfi <= ~MAH | mci; 
			nfj <= ~MAG | mch; 
			nfk <= MAF & mcg & ~MEH | ~MAF & ~mcg & ~MEH | ~MAF & mcg & MEH | ~MAF & mcg & ~MEH;
			nfl <= MAE & mcf & ~MEE | ~MAE & ~mcf & ~MEE | ~MAE & mcf & MEE | ~MAE & mcf & ~MEE;
			nfm <= MAD & mce & ~MEF | ~MAD & ~mce & ~MEF | ~MAD & mce & MEF | ~MAD & mce & ~MEF;
			nfn <= MAC & mcd & ~MED | ~MAC & ~mcd & ~MED | ~MAC & mcd & MED | ~MAC & mcd & ~MED;
			nfo <= MAB & mcc & ~MEB | ~MAB & ~mcc & ~MEB | ~MAB & mcc & MEB | ~MAB & mcc & ~MEB;
			nfp <= MAA & mcb & ~MEA | ~MAA & ~mcb & ~MEA | ~MAA & mcb & MEA | ~MAA & mcb & ~MEA;
			PAB <= NED; 
			PAC <= NED & ~nxb | NHE; 
			PAD <= NED & ~nxb & ~nxc | NHE & ~nxc | NIE; 
			PAE <= NED & ~nxb & ~nxc & ~nxd | NHE & ~nxc & ~nxd | NIE & ~nxd | NJE; 
			PAF <= NED & ~nxb & ~nxc & ~nxd & ~nxe | NHE & ~nxc & ~nxd & ~nxe | NIE & ~nxd & ~nxe | NJE & ~nxe & ~nxe | NKE; 
			PAG <= NHE & ~nxc & ~nxd & ~nxe & ~nxf | NIE & ~nxd & ~nxe & ~nxf | NJE & ~nxe & ~nxf | NKE & ~nxf & ~nxf | NLE; 
			PAH <= NIE & ~nxd & ~nxe & ~nxf & ~nxg | NJE & ~nxe & ~nxf & ~nxg | NKE & ~nxf & ~nxg | NLE & ~nxg & ~nxg | NME; 
			pai <= nxc | nxd | nxe | nxf | nxg; 
			pak <= ~NED | nxi | nxj | nxk | nxl; 
			PAL <= NHE; 
			PBA <= NAA; 
			PBB <= NAB; 
			PBC <= NAC; 
			PBD <= NAD; 
			PBE <= NAE; 
			PBF <= NAF & nee | ~NAF & ~nee; 
			PBG <= NAG & ~NHC | ~NAG & NHC; 
			PBH <= NAH & ~NHD | ~NAH & NHD; 
			PBI <= NAI; 
			PBJ <= NAJ & nei | ~NAJ & ~nei; 
			PBK <= NAK & ~NIC | ~NAK & NIC; 
			PBL <= NAL & ~NID | ~NAL & NID; 
			PBM <= NAM; 
			PBN <= NAN & nem | ~NAN & ~nem; 
			PBO <= NAO & ~NJC | ~NAO & NJC; 
			PBP <= NAP & ~NJD | ~NAP & NJD; 
			PCA <= NBA; 
			PCB <= NBB & nfa | ~NBB & ~nfa; 
			PCC <= NBC & ~NKC | ~NBC & NKC; 
			PCD <= NBD & ~NKD | ~NBD & NKD; 
			PCE <= NBE; 
			PCF <= NBF & nfe | ~NBF & ~nfe; 
			PCG <= NBG & ~NLC | ~NBG & NLC; 
			PCH <= NBH & ~NLD | ~NBH & NLD; 
			PCI <= NBI; 
			PCJ <= NBJ & nfi | ~NBJ & ~nfi; 
			PCK <= NBK & ~NMC | ~NBK & NMC; 
			PCL <= NBL & ~NMD | ~NBL & NMD; 
			PCM <= NBM; 
			PCN <= NBN & nfn | ~NBN & ~nfn; 
			PCO <= NBO & ~NNC | ~NBO & NNC; 
			PCP <= NBP & ~NND | ~NBP & NND; 
			PDE <= ~NAE; 
			PDF <= NAF & ~NAE | ~NAF & NAE; 
			PDG <= NAG & ~NPC | ~NAG & NPC; 
			PDH <= NAH & ~NPD | ~NAH & NPD; 
			PDI <= ~NAI; 
			PDJ <= NAJ & ~NAI | ~NAJ & NAI; 
			PDK <= NAK & ~NQC | ~NAK & NQC; 
			PDL <= NAL & ~NQD | ~NAL & NQD; 
			PDM <= ~NAM; 
			PDN <= NAN & ~NAM | ~NAN & NAM; 
			PDO <= NAO & ~NRC | ~NAO & NRC; 
			PDP <= NAP & ~NRD | ~NAP & NRD; 
			PEA <= ~NBA; 
			PEB <= NBB & ~NBA | ~NBB & NBA; 
			PEC <= NBC & ~NSC | ~NBC & NSC; 
			PED <= NBD & ~NSD | ~NBD & NSD; 
			PEE <= ~NBE; 
			PEF <= NBF & ~NBE | ~NBF & NBE; 
			PEG <= NBG & ~NTC | ~NBG & NTC; 
			PEH <= NBH & ~NTD | ~NBH & NTD; 
			PEI <= ~NBI; 
			PEJ <= NBJ & ~NBI | ~NBJ & NBI; 
			PEK <= NBK & ~NUC | ~NBK & NUC; 
			PEL <= NBL & ~NUD | ~NBL & NUD; 
			PEM <= ~NBM; 
			PEN <= NBN & ~NBM | ~NBN & NBM; 
			PEO <= NBO & ~NVC | ~NBO & NVC; 
			PEP <= NBP & ~NVD | ~NBP & NVD; 
			PFA <= PBA; 
			PFB <= PBB; 
			PFC <= PBC; 
			PFD <= PBD; 
			PFE <= PDE & PAB | PBE & ~PAB; 
			PFF <= PDF & PAB | PBF & ~PAB; 
			PFG <= PDG & PAB | PBG & ~PAB; 
			PFH <= PDH & PAB | PBH & ~PAB; 
			PFI <= PDI & PAC | PBI & ~PAC; 
			PFJ <= PDJ & PAC | PBJ & ~PAC; 
			PFK <= PDK & PAC | PBK & ~PAC; 
			PFL <= PDL & PAC | PBL & ~PAC; 
			PFM <= PDM & PAD | PBM & ~PAD; 
			PFN <= PDN & PAD | PBN & ~PAD; 
			PFO <= PDO & PAD | PBO & ~PAD; 
			PFP <= PDP & PAD | PBP & ~PAD; 
			PGA <= PEA & PAE | PCA & ~PAE; 
			PGB <= PEB & PAE | PCB & ~PAE; 
			PGC <= PEC & PAE | PCC & ~PAE; 
			PGD <= PED & PAE | PCD & ~PAE; 
			PGE <= PEE & PAF | PCE & ~PAF; 
			PGF <= PEF & PAF | PCF & ~PAF; 
			PGG <= PEG & PAF | PCG & ~PAF; 
			PGH <= PEH & PAF | PCH & ~PAF; 
			PGI <= PCI & ~PAG & pak | PEI & PAG | PEI & ~pak; 
			PGJ <= PCJ & ~PAG & pak | PEJ & PAG | PEJ & ~pak; 
			PGK <= PCK & ~PAG & pak | PEK & PAG | PEK & ~pak; 
			PGL <= PCL & ~PAG & pak | PEL & PAG | PEL & ~pak; 
			PGM <= PCM & ~PAH & ~PAM | PEM & PAH | PEM & PAM; 
			PGN <= PCN & ~PAH & ~PAM | PEN & PAH | PEN & PAM; 
			PGO <= PCO & ~PAH & ~PAM | PEO & PAH | PEO & PAM; 
			PGP <= PCP & ~PAH & ~PAM | PEP & PAH | PEP & PAM; 
			TFA <= QAI; 
			TFB <= QAI; 
			TFC <= QAI; 
			TFD <= QAI; 
			OAA <= PFA & TFA | ICA & ~TFA; 
			OAB <= PFB & TFA | ICB & ~TFA; 
			OAC <= PFC & TFA | ICC & ~TFA; 
			OAD <= PFD & TFA | ICD & ~TFA; 
			OAE <= PFE & TFA | ICE & ~TFA; 
			OAF <= PFF & TFA | ICF & ~TFA; 
			OAG <= PFG & TFA | ICG & ~TFA; 
			OAH <= PFH & TFA | ICH & ~TFA; 
			OAI <= PFI & TFB | ICI & ~TFB; 
			OAJ <= PFJ & TFB | ICJ & ~TFB; 
			OAK <= PFK & TFB | ICK & ~TFB; 
			OAL <= PFL & TFB | ICL & ~TFB; 
			OAM <= PFM & TFB | ICM & ~TFB; 
			OAN <= PFN & TFB | ICN & ~TFB; 
			OAO <= PFO & TFB | ICO & ~TFB; 
			OAP <= PFP & TFB | ICP & ~TFB; 
			OBA <= PGA & TFC | IDA & ~TFC; 
			OBB <= PGB & TFC | IDB & ~TFC; 
			OBC <= PGC & TFC | IDC & ~TFC; 
			OBD <= PGD & TFC | IDD & ~TFC; 
			OBE <= PGE & TFC | IDE & ~TFC; 
			OBF <= PGF & TFC | IDF & ~TFC; 
			OBG <= PGG & TFC | IDG & ~TFC; 
			OBH <= PGH & TFC | IDH & ~TFC; 
			OBI <= PGI & TFD | IDI & ~TFD; 
			OBJ <= PGJ & TFD | IDJ & ~TFD; 
			OBK <= PGK & TFD | IDK & ~TFD; 
			OBL <= PGL & TFD | IDL & ~TFD; 
			OBM <= PGM & TFD | IDM & ~TFD; 
			OBN <= PGN & TFD | IDN & ~TFD; 
			OBO <= PGO & TFD | IDO & ~TFD; 
			OBP <= PGP & TFD | IDP & ~TFD; 
			OEA <= IEA; 
			OEB <= IEB; 
			OEC <= IEC; 
			OED <= IED; 
			OEE <= IEE; 
			OEF <= IEF; 
			OFA <= IEA; 
			OFB <= IEB; 
			OFC <= IEC; 
			OFD <= IED; 
			OFE <= IEE; 
			OFF <= IEF; 
			OJA <= IFA; 
			OJB <= IFB; 
			OJC <= IFC; 
			OJD <= IFD; 
			OJE <= IFE; 
			OJF <= IFF; 
			OJG <= IFG; 
			OJH <= IGA; 
			OJI <= IGB; 
			OJJ <= IGC; 
			OJK <= IGD; 
			OJL <= IGE; 
			OJM <= IGF; 
			OLA <= IFA; 
			OLB <= IFB; 
			OLC <= IFC; 
			OLD <= IFD; 
			OLE <= IFE; 
			OLF <= IFF; 
			OLG <= IFG; 
			OLH <= IGA; 
			OLI <= IGB; 
			OLJ <= IGC; 
			OLK <= IGD; 
			OLL <= IGE; 
			OLM <= IGF; 
			ONA <= IFA; 
			ONB <= IFB; 
			ONC <= IFC; 
			OND <= IFD; 
			ONE <= IFE; 
			ONF <= IFF; 
			ONG <= IFG; 
			ONH <= IGA; 
			ONI <= IGB; 
			ONJ <= IGC; 
			ONK <= IGD; 
			ONL <= IGE; 
			ONM <= IGF; 
			OPA <= IFA; 
			OPB <= IFB; 
			OPC <= IFC; 
			OPD <= IFD; 
			OPE <= IFE; 
			OPF <= IFF; 
			OPG <= IFG; 
			OPH <= IGA; 
			OPI <= IGB; 
			OPJ <= IGC; 
			OPK <= IGD; 
			OPL <= IGE; 
			OPM <= IGF;			
		end 
endmodule
