module fb( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IAR, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBM, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFF, 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IJA, 
 IJB, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 OEA, 
 OEB, 
 OFA, 
 OFB, 
 OGA, 
 OGB, 
 OHA, 
 OHB, 
 OIA, 
 OJA, 
OJB ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IAR; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBM; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFF; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IJA; 
 input IJB; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output OEA; 
 output OEB; 
 output OFA; 
 output OFB; 
 output OGA; 
 output OGB; 
 output OHA; 
 output OHB; 
 output OIA; 
 output OJA; 
 output OJB; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  AAQ ;
reg  aar ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  baa ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FBA ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FDA ;
reg  FDB ;
reg  FDC ;
reg  FDD ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FFA ;
reg  FFB ;
reg  FFC ;
reg  FFD ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FHA ;
reg  FHB ;
reg  FHC ;
reg  FHD ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FJA ;
reg  FJB ;
reg  FJC ;
reg  FJD ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FLA ;
reg  FLB ;
reg  FLC ;
reg  FLD ;
reg  gba ;
reg  gca ;
reg  gda ;
reg  GEA ;
reg  GEB ;
reg  GEC ;
reg  GED ;
reg  gfa ;
reg  gga ;
reg  gha ;
reg  GIA ;
reg  GIB ;
reg  GIC ;
reg  GID ;
reg  gja ;
reg  gka ;
reg  gla ;
reg  GMA ;
reg  GMB ;
reg  GMC ;
reg  GMD ;
reg  haa ;
reg  hab ;
reg  hac ;
reg  had ;
reg  hae ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hce ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  KCD ;
reg  KCE ;
reg  KCF ;
reg  KCG ;
reg  KCH ;
reg  KDA ;
reg  KDB ;
reg  KDC ;
reg  KDD ;
reg  KDE ;
reg  KDF ;
reg  KDG ;
reg  KDH ;
reg  KEA ;
reg  KEB ;
reg  KEC ;
reg  KED ;
reg  KEE ;
reg  KEF ;
reg  KEG ;
reg  KEH ;
reg  KFA ;
reg  KFB ;
reg  KFC ;
reg  KFD ;
reg  KFE ;
reg  KFF ;
reg  KFG ;
reg  KFH ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  KGD ;
reg  KGE ;
reg  KGF ;
reg  KGG ;
reg  KGH ;
reg  KHA ;
reg  KHB ;
reg  KHC ;
reg  KHD ;
reg  KHE ;
reg  KHF ;
reg  KHG ;
reg  KHH ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  KID ;
reg  KIE ;
reg  KIF ;
reg  KIG ;
reg  KIH ;
reg  KJA ;
reg  KJB ;
reg  KJC ;
reg  KJD ;
reg  KJE ;
reg  KJF ;
reg  KJG ;
reg  KJH ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  KKD ;
reg  KKE ;
reg  KKF ;
reg  KKG ;
reg  KKH ;
reg  KLA ;
reg  KLB ;
reg  KLC ;
reg  KLD ;
reg  KLE ;
reg  KLF ;
reg  KLG ;
reg  KLH ;
reg  naa ;
reg  nab ;
reg  nac ;
reg  nad ;
reg  nae ;
reg  naf ;
reg  nag ;
reg  nah ;
reg  nai ;
reg  naj ;
reg  nak ;
reg  nal ;
reg  nba ;
reg  nbb ;
reg  nbc ;
reg  nbd ;
reg  nbe ;
reg  nbf ;
reg  nbg ;
reg  nbh ;
reg  nbi ;
reg  nbj ;
reg  nbk ;
reg  nbl ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ode ;
reg  OEA ;
reg  OEB ;
reg  OFA ;
reg  OFB ;
reg  OGA ;
reg  OGB ;
reg  oha ;
reg  OHB ;
reg  OIA ;
reg  oja ;
reg  ojb ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  qbf ;
reg  qbg ;
reg  qbh ;
reg  QCA ;
reg  QDA ;
reg  QDB ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  QFA ;
reg  QFB ;
reg  qga ;
reg  UAA ;
reg  UAB ;
reg  UBA ;
reg  UBB ;
reg  UCA ;
reg  UCB ;
reg  UDA ;
reg  UDB ;
reg  UEA ;
reg  UEB ;
reg  UFA ;
reg  UFB ;
reg  UGA ;
reg  UGB ;
reg  UHA ;
reg  UHB ;
reg  UIA ;
reg  UIB ;
reg  UJA ;
reg  UJB ;
reg  UKA ;
reg  UKB ;
reg  ULA ;
reg  ULB ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aaq ;
wire  AAR ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  BAA ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  caf ;
wire  CAF ;
wire  cag ;
wire  CAG ;
wire  cah ;
wire  CAH ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cbe ;
wire  CBE ;
wire  cbf ;
wire  CBF ;
wire  cbg ;
wire  CBG ;
wire  cbh ;
wire  CBH ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cce ;
wire  CCE ;
wire  ccf ;
wire  CCF ;
wire  ccg ;
wire  CCG ;
wire  cch ;
wire  CCH ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cde ;
wire  CDE ;
wire  cdf ;
wire  CDF ;
wire  cdg ;
wire  CDG ;
wire  cdh ;
wire  CDH ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cee ;
wire  CEE ;
wire  cef ;
wire  CEF ;
wire  ceg ;
wire  CEG ;
wire  ceh ;
wire  CEH ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cfe ;
wire  CFE ;
wire  cff ;
wire  CFF ;
wire  cfg ;
wire  CFG ;
wire  cfh ;
wire  CFH ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cge ;
wire  CGE ;
wire  cgf ;
wire  CGF ;
wire  cgg ;
wire  CGG ;
wire  cgh ;
wire  CGH ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  che ;
wire  CHE ;
wire  chf ;
wire  CHF ;
wire  chg ;
wire  CHG ;
wire  chh ;
wire  CHH ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cie ;
wire  CIE ;
wire  cif ;
wire  CIF ;
wire  cig ;
wire  CIG ;
wire  cih ;
wire  CIH ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cje ;
wire  CJE ;
wire  cjf ;
wire  CJF ;
wire  cjg ;
wire  CJG ;
wire  cjh ;
wire  CJH ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cke ;
wire  CKE ;
wire  ckf ;
wire  CKF ;
wire  ckg ;
wire  CKG ;
wire  ckh ;
wire  CKH ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cle ;
wire  CLE ;
wire  clf ;
wire  CLF ;
wire  clg ;
wire  CLG ;
wire  clh ;
wire  CLH ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  eee ;
wire  EEE ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  efe ;
wire  EFE ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  ege ;
wire  EGE ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  ehe ;
wire  EHE ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eic ;
wire  EIC ;
wire  eid ;
wire  EID ;
wire  eie ;
wire  EIE ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eje ;
wire  EJE ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ekd ;
wire  EKD ;
wire  eke ;
wire  EKE ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ele ;
wire  ELE ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fba ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fda ;
wire  fdb ;
wire  fdc ;
wire  fdd ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  ffa ;
wire  ffb ;
wire  ffc ;
wire  ffd ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fha ;
wire  fhb ;
wire  fhc ;
wire  fhd ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fja ;
wire  fjb ;
wire  fjc ;
wire  fjd ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fla ;
wire  flb ;
wire  flc ;
wire  fld ;
wire  GBA ;
wire  GCA ;
wire  GDA ;
wire  gea ;
wire  geb ;
wire  gec ;
wire  ged ;
wire  GFA ;
wire  GGA ;
wire  GHA ;
wire  gia ;
wire  gib ;
wire  gic ;
wire  gid ;
wire  GJA ;
wire  GKA ;
wire  GLA ;
wire  gma ;
wire  gmb ;
wire  gmc ;
wire  gmd ;
wire  HAA ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  HAE ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HCE ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iar ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibm ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iff ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  ija ;
wire  ijb ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  kcd ;
wire  kce ;
wire  kcf ;
wire  kcg ;
wire  kch ;
wire  kda ;
wire  kdb ;
wire  kdc ;
wire  kdd ;
wire  kde ;
wire  kdf ;
wire  kdg ;
wire  kdh ;
wire  kea ;
wire  keb ;
wire  kec ;
wire  ked ;
wire  kee ;
wire  kef ;
wire  keg ;
wire  keh ;
wire  kfa ;
wire  kfb ;
wire  kfc ;
wire  kfd ;
wire  kfe ;
wire  kff ;
wire  kfg ;
wire  kfh ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  kgd ;
wire  kge ;
wire  kgf ;
wire  kgg ;
wire  kgh ;
wire  kha ;
wire  khb ;
wire  khc ;
wire  khd ;
wire  khe ;
wire  khf ;
wire  khg ;
wire  khh ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  kid ;
wire  kie ;
wire  kif ;
wire  kig ;
wire  kih ;
wire  kja ;
wire  kjb ;
wire  kjc ;
wire  kjd ;
wire  kje ;
wire  kjf ;
wire  kjg ;
wire  kjh ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  kkd ;
wire  kke ;
wire  kkf ;
wire  kkg ;
wire  kkh ;
wire  kla ;
wire  klb ;
wire  klc ;
wire  kld ;
wire  kle ;
wire  klf ;
wire  klg ;
wire  klh ;
wire  maa ;
wire  MAA ;
wire  mab ;
wire  MAB ;
wire  mac ;
wire  MAC ;
wire  mad ;
wire  MAD ;
wire  mae ;
wire  MAE ;
wire  maf ;
wire  MAF ;
wire  mag ;
wire  MAG ;
wire  mah ;
wire  MAH ;
wire  mai ;
wire  MAI ;
wire  maj ;
wire  MAJ ;
wire  mak ;
wire  MAK ;
wire  mal ;
wire  MAL ;
wire  mba ;
wire  MBA ;
wire  mbb ;
wire  MBB ;
wire  mbc ;
wire  MBC ;
wire  mbd ;
wire  MBD ;
wire  mbe ;
wire  MBE ;
wire  mbf ;
wire  MBF ;
wire  mbg ;
wire  MBG ;
wire  mbh ;
wire  MBH ;
wire  mbi ;
wire  MBI ;
wire  mbj ;
wire  MBJ ;
wire  mbk ;
wire  MBK ;
wire  mbl ;
wire  MBL ;
wire  mca ;
wire  MCA ;
wire  mcb ;
wire  MCB ;
wire  mcc ;
wire  MCC ;
wire  mcd ;
wire  MCD ;
wire  mce ;
wire  MCE ;
wire  mcf ;
wire  MCF ;
wire  mcg ;
wire  MCG ;
wire  mch ;
wire  MCH ;
wire  mci ;
wire  MCI ;
wire  mcj ;
wire  MCJ ;
wire  mck ;
wire  MCK ;
wire  mcl ;
wire  MCL ;
wire  mda ;
wire  MDA ;
wire  mdb ;
wire  MDB ;
wire  mdc ;
wire  MDC ;
wire  mdd ;
wire  MDD ;
wire  mde ;
wire  MDE ;
wire  mdf ;
wire  MDF ;
wire  mdg ;
wire  MDG ;
wire  mdh ;
wire  MDH ;
wire  mdi ;
wire  MDI ;
wire  mdj ;
wire  MDJ ;
wire  mdk ;
wire  MDK ;
wire  mdl ;
wire  MDL ;
wire  NAA ;
wire  NAB ;
wire  NAC ;
wire  NAD ;
wire  NAE ;
wire  NAF ;
wire  NAG ;
wire  NAH ;
wire  NAI ;
wire  NAJ ;
wire  NAK ;
wire  NAL ;
wire  NBA ;
wire  NBB ;
wire  NBC ;
wire  NBD ;
wire  NBE ;
wire  NBF ;
wire  NBG ;
wire  NBH ;
wire  NBI ;
wire  NBJ ;
wire  NBK ;
wire  NBL ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ODE ;
wire  oea ;
wire  oeb ;
wire  ofa ;
wire  ofb ;
wire  oga ;
wire  ogb ;
wire  OHA ;
wire  ohb ;
wire  oia ;
wire  OJA ;
wire  OJB ;
wire  paa ;
wire  PAA ;
wire  pab ;
wire  PAB ;
wire  pac ;
wire  PAC ;
wire  pba ;
wire  PBA ;
wire  pbb ;
wire  PBB ;
wire  pbc ;
wire  PBC ;
wire  pbd ;
wire  PBD ;
wire  pca ;
wire  PCA ;
wire  pcb ;
wire  PCB ;
wire  pcc ;
wire  PCC ;
wire  pcd ;
wire  PCD ;
wire  pda ;
wire  PDA ;
wire  pdb ;
wire  PDB ;
wire  pdc ;
wire  PDC ;
wire  pdd ;
wire  PDD ;
wire  peb ;
wire  PEB ;
wire  pec ;
wire  PEC ;
wire  pfb ;
wire  PFB ;
wire  pfc ;
wire  PFC ;
wire  pgb ;
wire  PGB ;
wire  pgc ;
wire  PGC ;
wire  phb ;
wire  PHB ;
wire  phc ;
wire  PHC ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  QBF ;
wire  QBG ;
wire  QBH ;
wire  qca ;
wire  qda ;
wire  qdb ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  qfa ;
wire  qfb ;
wire  QGA ;
wire  raa ;
wire  RAA ;
wire  rab ;
wire  RAB ;
wire  rba ;
wire  RBA ;
wire  rbb ;
wire  RBB ;
wire  rca ;
wire  RCA ;
wire  rcb ;
wire  RCB ;
wire  rda ;
wire  RDA ;
wire  rdb ;
wire  RDB ;
wire  rea ;
wire  REA ;
wire  reb ;
wire  REB ;
wire  rfa ;
wire  RFA ;
wire  rfb ;
wire  RFB ;
wire  rga ;
wire  RGA ;
wire  rgb ;
wire  RGB ;
wire  rha ;
wire  RHA ;
wire  rhb ;
wire  RHB ;
wire  ria ;
wire  RIA ;
wire  rib ;
wire  RIB ;
wire  rja ;
wire  RJA ;
wire  rjb ;
wire  RJB ;
wire  rka ;
wire  RKA ;
wire  rkb ;
wire  RKB ;
wire  rla ;
wire  RLA ;
wire  rlb ;
wire  RLB ;
wire  saa ;
wire  SAA ;
wire  sab ;
wire  SAB ;
wire  sac ;
wire  SAC ;
wire  sad ;
wire  SAD ;
wire  sba ;
wire  SBA ;
wire  sbb ;
wire  SBB ;
wire  sbc ;
wire  SBC ;
wire  sbd ;
wire  SBD ;
wire  sca ;
wire  SCA ;
wire  scb ;
wire  SCB ;
wire  scc ;
wire  SCC ;
wire  scd ;
wire  SCD ;
wire  sda ;
wire  SDA ;
wire  sdb ;
wire  SDB ;
wire  sdc ;
wire  SDC ;
wire  sdd ;
wire  SDD ;
wire  sea ;
wire  SEA ;
wire  seb ;
wire  SEB ;
wire  sec ;
wire  SEC ;
wire  sed ;
wire  SED ;
wire  sfa ;
wire  SFA ;
wire  sfb ;
wire  SFB ;
wire  sfc ;
wire  SFC ;
wire  sfd ;
wire  SFD ;
wire  sga ;
wire  SGA ;
wire  sgb ;
wire  SGB ;
wire  sgc ;
wire  SGC ;
wire  sgd ;
wire  SGD ;
wire  sha ;
wire  SHA ;
wire  shb ;
wire  SHB ;
wire  shc ;
wire  SHC ;
wire  shd ;
wire  SHD ;
wire  sia ;
wire  SIA ;
wire  sib ;
wire  SIB ;
wire  sic ;
wire  SIC ;
wire  sid ;
wire  SID ;
wire  sja ;
wire  SJA ;
wire  sjb ;
wire  SJB ;
wire  sjc ;
wire  SJC ;
wire  sjd ;
wire  SJD ;
wire  ska ;
wire  SKA ;
wire  skb ;
wire  SKB ;
wire  skc ;
wire  SKC ;
wire  skd ;
wire  SKD ;
wire  sla ;
wire  SLA ;
wire  slb ;
wire  SLB ;
wire  slc ;
wire  SLC ;
wire  sld ;
wire  SLD ;
wire  uaa ;
wire  uab ;
wire  uba ;
wire  ubb ;
wire  uca ;
wire  ucb ;
wire  uda ;
wire  udb ;
wire  uea ;
wire  ueb ;
wire  ufa ;
wire  ufb ;
wire  uga ;
wire  ugb ;
wire  uha ;
wire  uhb ;
wire  uia ;
wire  uib ;
wire  uja ;
wire  ujb ;
wire  uka ;
wire  ukb ;
wire  ula ;
wire  ulb ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign jam =  ZZO & ged & gic & gmb  |  ZZI & ged & gic & gmb  |  hbd & gic & gmb  |  hcd & gmb  ; 
assign JAM = ~jam;  //complement 
assign gid = ~GID;  //complement 
assign OHA = ~oha;  //complement 
assign QGA = ~qga;  //complement 
assign JBC =  ZZO & gec & gid & gmd & QAG  |  ZZI & gec & gid & gmd & QAG  |  hbe & gid & gmd & QAG  |  hce & gmd & QAG  |  ZZO & QAG  |  QCA  ; 
assign jbc = ~JBC;  //complement 
assign GCA = ~gca;  //complement 
assign ohb = ~OHB;  //complement 
assign RKA =  UKA & qbh & qbh  |  UKB & QBH & QBH  ; 
assign rka = ~RKA;  //complement 
assign RKB =  fkd & fkc & qbh  |  FKD & FKC & QBH  ; 
assign rkb = ~RKB;  //complement 
assign oca = ~OCA;  //complement 
assign ocb = ~OCB;  //complement 
assign occ = ~OCC;  //complement 
assign RIA =  UIA & qbh & qbh  |  UIB & QBH & QBH  ; 
assign ria = ~RIA;  //complement 
assign RIB =  fid & fic & qbh  |  FID & FIC & QBH  ; 
assign rib = ~RIB;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign ocd = ~OCD;  //complement 
assign QBE = ~qbe;  //complement 
assign QBF = ~qbf;  //complement 
assign QBG = ~qbg;  //complement 
assign QBH = ~qbh;  //complement 
assign RGB =  ffd & fgc & qbh  |  FGD & FGC & QBH  ; 
assign rgb = ~RGB;  //complement 
assign RGA =  UGA & qbh & qbh  |  UGB & QBH & QBH  ; 
assign rga = ~RGA;  //complement 
assign ODE = ~ode;  //complement 
assign obk = ~OBK;  //complement 
assign obl = ~OBL;  //complement 
assign oci = ~OCI;  //complement 
assign QBA = ~qba;  //complement 
assign QBB = ~qbb;  //complement 
assign QBC = ~qbc;  //complement 
assign QBD = ~qbd;  //complement 
assign ofa = ~OFA;  //complement 
assign oga = ~OGA;  //complement 
assign ocj = ~OCJ;  //complement 
assign ock = ~OCK;  //complement 
assign ocl = ~OCL;  //complement 
assign HAA = ~haa;  //complement 
assign HAB = ~hab;  //complement 
assign oea = ~OEA;  //complement 
assign odc = ~ODC;  //complement 
assign ocm = ~OCM;  //complement 
assign ocn = ~OCN;  //complement 
assign oco = ~OCO;  //complement 
assign RHA =  UHA & qbg & qbg  |  UHB & QBG & QBG  ; 
assign rha = ~RHA;  //complement 
assign RHB =  fhd & fhc & qbg  |  FHD & FHC & QBG  ; 
assign rhb = ~RHB;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign ocp = ~OCP;  //complement 
assign RJA =  UJA & qbg & qbg  |  UJB & QBG & QBG  ; 
assign rja = ~RJA;  //complement 
assign RJB =  fjd & fjc & qbg  |  FJD & FJC & QBG  ; 
assign rjb = ~RJB;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign oce = ~OCE;  //complement 
assign RLA =  ULA & qbg & qbg  |  ULB & QBG & QBG  ; 
assign rla = ~RLA;  //complement 
assign RLB =  fld & flc & qbg  |  FLD & FLC & QBG  ; 
assign rlb = ~RLB;  //complement 
assign ocf = ~OCF;  //complement 
assign ocg = ~OCG;  //complement 
assign och = ~OCH;  //complement 
assign qab = ~QAB;  //complement 
assign qca = ~QCA;  //complement 
assign qfa = ~QFA;  //complement 
assign qaa = ~QAA;  //complement 
assign JBB =  ZZO & ged & gic & gmb & QAG  |  ZZI & ged & gic & gmb & QAG  |  hbd & gic & gmb & QAG  |  hcd & gmb & QAG  |  ZZO & QAG  |  QCA  ; 
assign jbb = ~JBB;  //complement 
assign gic = ~GIC;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign JBA =  ZZO & gec & gid & gmd & QAG  |  ZZI & gec & gid & gmd & QAG  |  hbe & gid & gmd & QAG  |  hce & gmd & QAG  |  ZZO & QAG  |  QCA  ; 
assign jba = ~JBA;  //complement 
assign gec = ~GEC;  //complement 
assign REA =  UEA & qbf & qbf  |  UEB & QBF & QBF  ; 
assign rea = ~REA;  //complement 
assign REB =  fed & fec & qbf  |  FED & FEC & QBF  ; 
assign reb = ~REB;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign oak = ~OAK;  //complement 
assign RCA =  UCA & qbf & qbf  |  UCB & QBF & QBF  ; 
assign rca = ~RCA;  //complement 
assign RCB =  fcd & fcc & qbf  |  FCD & FCC & QBF  ; 
assign rcb = ~RCB;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign oal = ~OAL;  //complement 
assign RAA =  UAA & qbf & qbf  |  UAB & QBF & QBF  ; 
assign raa = ~RAA;  //complement 
assign RAB =  fad & fac & qbf  |  FAD & FAC & QBF  ; 
assign rab = ~RAB;  //complement 
assign oac = ~OAC;  //complement 
assign oad = ~OAD;  //complement 
assign oba = ~OBA;  //complement 
assign HBA = ~hba;  //complement 
assign HBB = ~hbb;  //complement 
assign ofb = ~OFB;  //complement 
assign ogb = ~OGB;  //complement 
assign obb = ~OBB;  //complement 
assign obc = ~OBC;  //complement 
assign obd = ~OBD;  //complement 
assign HAC = ~hac;  //complement 
assign oeb = ~OEB;  //complement 
assign odd = ~ODD;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign obg = ~OBG;  //complement 
assign qfb = ~QFB;  //complement 
assign OJB = ~ojb;  //complement 
assign RBA =  UBA & qbe & qbe  |  UBB & QBE & QBE  ; 
assign rba = ~RBA;  //complement 
assign RBB =  fbd & fbc & qbe  |  FBD & FBC & QBE  ; 
assign rbb = ~RBB;  //complement 
assign OJA = ~oja;  //complement 
assign QEA = ~qea;  //complement 
assign QEB = ~qeb;  //complement 
assign QEC = ~qec;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign obh = ~OBH;  //complement 
assign RDA =  UDA & qbe & qbe  |  UDB & QBE & QBE  ; 
assign rda = ~RDA;  //complement 
assign RDB =  fdd & fdc & qbe  |  FDD & FDC & QBE  ; 
assign rdb = ~RDB;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign oam = ~OAM;  //complement 
assign RFA =  UFA & qbe & qbe  |  UFB & QBE & QBE  ; 
assign rfa = ~RFA;  //complement 
assign RFB =  ffd & ffc & qbe  |  FFD & FFC & QBE  ; 
assign rfb = ~RFB;  //complement 
assign oan = ~OAN;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign MAK =  kka & kkb & kkc & kkd  ; 
assign mak = ~MAK;  //complement  
assign MBK =  kke & kkf & kkg & kkh  ; 
assign mbk = ~MBK;  //complement 
assign MAL =  kla & klb & klc & kld  ; 
assign mal = ~MAL;  //complement  
assign MBL =  kle & klf & klg & klh  ; 
assign mbl = ~MBL;  //complement 
assign MCK =  KKA & KKB & KKC & KKD  ; 
assign mck = ~MCK;  //complement  
assign MDK =  KKE & KKF & KKG & KKH  ; 
assign mdk = ~MDK;  //complement 
assign fka = ~FKA;  //complement 
assign fkb = ~FKB;  //complement 
assign kkb = ~KKB;  //complement 
assign kkf = ~KKF;  //complement 
assign ska =  kkc & KKB  |  KKD  ; 
assign SKA = ~ska;  //complement 
assign skb =  KKC & kkb  |  kkd  ; 
assign SKB = ~skb;  //complement 
assign fkc = ~FKC;  //complement 
assign fkd = ~FKD;  //complement 
assign kkd = ~KKD;  //complement 
assign kkh = ~KKH;  //complement 
assign skc =  kkg & KKF  |  KKH  ; 
assign SKC = ~skc;  //complement 
assign skd =  KKG & kkf  |  kkh  ; 
assign SKD = ~skd;  //complement 
assign fla = ~FLA;  //complement 
assign flb = ~FLB;  //complement 
assign NAK = ~nak;  //complement 
assign NBK = ~nbk;  //complement 
assign uka = ~UKA;  //complement 
assign ukb = ~UKB;  //complement 
assign pda =  naj & nbj  |  nak & nbk  |  nal & nbl  ; 
assign PDA = ~pda;  //complement 
assign pac =  nai & nbi  |  naj & nbj  |  nak & nbk  |  nal & nbl  ; 
assign PAC = ~pac;  //complement 
assign pec =  nai & nbi  |  naj & nbj  |  nak & nbk  |  nal & nbl  ; 
assign PEC = ~pec; //complement 
assign gib = ~GIB;  //complement 
assign pdc =  nal & nbl  |  NAK  |  NBK  ; 
assign PDC = ~pdc;  //complement 
assign phc =  nal & nbl  |  NAK  |  NBK  ; 
assign PHC = ~phc; //complement 
assign pdb =  NAJ  |  NBJ  |  nak & nbk  |  nal & nbl  ; 
assign PDB = ~pdb;  //complement 
assign phb =  NAJ  |  NBJ  |  nak & nbk  |  nal & nbl  ; 
assign PHB = ~phb; //complement 
assign ged = ~GED;  //complement 
assign slc =  klg & KLF  |  KLH  ; 
assign SLC = ~slc;  //complement 
assign sld =  KLG & klf  |  klh  ; 
assign SLD = ~sld;  //complement 
assign NAL = ~nal;  //complement 
assign NBL = ~nbl;  //complement 
assign ula = ~ULA;  //complement 
assign ulb = ~ULB;  //complement 
assign sla =  klc & KLB  |  KLD  ; 
assign SLA = ~sla;  //complement 
assign slb =  KLC & klb  |  kld  ; 
assign SLB = ~slb;  //complement 
assign klb = ~KLB;  //complement 
assign klf = ~KLF;  //complement 
assign MCL =  KLA & KLB & KLC & KLD  ; 
assign mcl = ~MCL;  //complement  
assign MDL =  KLE & KLF & KLG & KLH  ; 
assign mdl = ~MDL;  //complement 
assign flc = ~FLC;  //complement 
assign fld = ~FLD;  //complement 
assign kld = ~KLD;  //complement 
assign klh = ~KLH;  //complement 
assign kka = ~KKA;  //complement 
assign kke = ~KKE;  //complement 
assign ckb =  bci  ; 
assign CKB = ~ckb;  //complement 
assign ckc =  bcj & bci  |  aci  ; 
assign CKC = ~ckc;  //complement 
assign aci = ~ACI;  //complement 
assign bci = ~BCI;  //complement 
assign kkc = ~KKC;  //complement 
assign kkg = ~KKG;  //complement 
assign CKF =  ACI  ; 
assign ckf = ~CKF;  //complement 
assign CKG =  ACJ & ACI  |  BCJ  ; 
assign ckg = ~CKG;  //complement 
assign ckd =  bci & bcj & bck  |  acj & bck  |  ack  ; 
assign CKD = ~ckd;  //complement 
assign acj = ~ACJ;  //complement 
assign bcj = ~BCJ;  //complement 
assign JAK =  GMA & HAD & QAF & HBD & HCB  |  ZZO & QAF & HBD & HCB  |  GEC & HBD & HCB  |  GEC & HCB  |  GKA  ; 
assign jak = ~JAK;  //complement 
assign CKH =  ACI & ACJ & ACK  |  BCJ & ACK  |  BCK  ; 
assign ckh = ~CKH;  //complement 
assign cke =  bci & bcj & bck & bcl  |  acj & bck & bcl  |  ack & bcl  |  acl  ; 
assign CKE = ~cke;  //complement 
assign ack = ~ACK;  //complement 
assign bck = ~BCK;  //complement 
assign HBD = ~hbd;  //complement 
assign HBE = ~hbe;  //complement 
assign EKD =  ACL & bcl  ; 
assign ekd = ~EKD;  //complement  
assign EKE =  ACI & ACJ & ACK & ACL  ; 
assign eke = ~EKE;  //complement 
assign EKA =  ACI & bci  ; 
assign eka = ~EKA;  //complement 
assign EKB =  ACJ & bcj  ; 
assign ekb = ~EKB;  //complement 
assign EKC =  ACK & bck  ; 
assign ekc = ~EKC;  //complement 
assign acl = ~ACL;  //complement 
assign bcl = ~BCL;  //complement 
assign HAD = ~had;  //complement 
assign HAE = ~hae;  //complement 
assign ELD =  ACP & bcp  ; 
assign eld = ~ELD;  //complement  
assign ELE =  ACM & ACN & ACO & ACP  ; 
assign ele = ~ELE;  //complement 
assign ELA =  ACM & bcm  ; 
assign ela = ~ELA;  //complement 
assign ELB =  ACN & bcn  ; 
assign elb = ~ELB;  //complement 
assign ELC =  ACO & bco  ; 
assign elc = ~ELC;  //complement 
assign acm = ~ACM;  //complement 
assign bcm = ~BCM;  //complement 
assign JAL =  GMD & HAE & QAE & HBE & HCC  |  ZZO & QAE & HBE & HCC  |  GED & HBE & HCC  |  GIB & HCC  |  GLA  ; 
assign jal = ~JAL;  //complement 
assign CLF =  ACM  ; 
assign clf = ~CLF;  //complement 
assign CLG =  ACN & ACM  |  BCN  ; 
assign clg = ~CLG;  //complement 
assign cle =  bcm & bcn & bco & bcp  |  acn & bco & bcp  |  aco & bcp  |  acp  ; 
assign CLE = ~cle;  //complement 
assign acn = ~ACN;  //complement 
assign bcn = ~BCN;  //complement 
assign kla = ~KLA;  //complement 
assign kle = ~KLE;  //complement 
assign CLH =  ACM & ACN & ACO  |  BCN & ACO  |  BCO  ; 
assign clh = ~CLH;  //complement 
assign cld =  bcm & bcn & bco  |  acn & bco  |  aco  ; 
assign CLD = ~cld;  //complement 
assign aco = ~ACO;  //complement 
assign bco = ~BCO;  //complement 
assign klc = ~KLC;  //complement 
assign klg = ~KLG;  //complement 
assign clb =  bcm  ; 
assign CLB = ~clb;  //complement 
assign clc =  bcn & bcm  |  acn  ; 
assign CLC = ~clc;  //complement 
assign acp = ~ACP;  //complement 
assign bcp = ~BCP;  //complement 
assign MAJ =  kja & kjb & kjc & kjd  ; 
assign maj = ~MAJ;  //complement  
assign MBJ =  kje & kjf & kjg & kjh  ; 
assign mbj = ~MBJ;  //complement 
assign MAI =  kia & kib & kic & kid  ; 
assign mai = ~MAI;  //complement  
assign MBI =  kie & kif & kig & kih  ; 
assign mbi = ~MBI;  //complement 
assign MCI =  KIA & KIB & KIC & KID  ; 
assign mci = ~MCI;  //complement  
assign MDI =  KIE & KIF & KIG & KIH  ; 
assign mdi = ~MDI;  //complement 
assign fia = ~FIA;  //complement 
assign fib = ~FIB;  //complement 
assign kib = ~KIB;  //complement 
assign kif = ~KIF;  //complement 
assign sia =  kic & KIB  |  KID  ; 
assign SIA = ~sia;  //complement 
assign sib =  KIC & kib  |  kid  ; 
assign SIB = ~sib;  //complement 
assign fic = ~FIC;  //complement 
assign kid = ~KID;  //complement 
assign kih = ~KIH;  //complement 
assign sic =  kig & KIF  |  KIH  ; 
assign SIC = ~sic;  //complement 
assign sid =  KIG & kif  |  kih  ; 
assign SID = ~sid;  //complement 
assign fja = ~FJA;  //complement 
assign fjb = ~FJB;  //complement 
assign NAI = ~nai;  //complement 
assign NBI = ~nbi;  //complement 
assign uia = ~UIA;  //complement 
assign uib = ~UIB;  //complement 
assign gia = ~GIA;  //complement 
assign kjb = ~KJB;  //complement 
assign kjf = ~KJF;  //complement 
assign pdd =  NAL  |  NBL  ; 
assign PDD = ~pdd;  //complement 
assign geb = ~GEB;  //complement 
assign sjc =  kjg & KJF  |  KJH  ; 
assign SJC = ~sjc;  //complement 
assign sjd =  KJG & kjf  |  kjh  ; 
assign SJD = ~sjd;  //complement 
assign NAJ = ~naj;  //complement 
assign NBJ = ~nbj;  //complement 
assign uja = ~UJA;  //complement 
assign ujb = ~UJB;  //complement 
assign sjb =  KJC & kjb  |  kid  ; 
assign SJB = ~sjb;  //complement 
assign fjc = ~FJC;  //complement 
assign fjd = ~FJD;  //complement 
assign MCJ =  KJA & KJB & KJC & KJD  ; 
assign mcj = ~MCJ;  //complement  
assign MDJ =  KJE & KJF & KJG & KJH  ; 
assign mdj = ~MDJ;  //complement 
assign pcd =  MAH  |  NBH  ; 
assign PCD = ~pcd;  //complement 
assign kjd = ~KJD;  //complement 
assign kjh = ~KJH;  //complement 
assign kia = ~KIA;  //complement 
assign kie = ~KIE;  //complement 
assign cib =  bca  ; 
assign CIB = ~cib;  //complement 
assign cic =  bcb & bca  |  acb  ; 
assign CIC = ~cic;  //complement 
assign aca = ~ACA;  //complement 
assign bca = ~BCA;  //complement 
assign kic = ~KIC;  //complement 
assign kig = ~KIG;  //complement 
assign CIF =  ACA  ; 
assign cif = ~CIF;  //complement 
assign CIG =  ACB & ACA  |  BCB  ; 
assign cig = ~CIG;  //complement 
assign cid =  bca & bcb & bcc  |  acb & bcc  |  acc  ; 
assign CID = ~cid;  //complement 
assign acb = ~ACB;  //complement 
assign bcb = ~BCB;  //complement 
assign JAI =  ZZO & QAF & HAD & HBD  |  GMA & QAF & HAD & HBD  |  ZZO & HAD & HBD  |  GEC & HBD  |  GID  ; 
assign jai = ~JAI;  //complement 
assign CIH =  ACA & ACB & ACC  |  BCB & ACC  |  BCC  ; 
assign cih = ~CIH;  //complement 
assign cie =  bca & bcb & bcc & bcd  |  acb & bcc & bcd  |  acc & bcd  |  acd  ; 
assign CIE = ~cie;  //complement 
assign acc = ~ACC;  //complement 
assign bcc = ~BCC;  //complement 
assign HBC = ~hbc;  //complement 
assign HCC = ~hcc;  //complement 
assign EID =  ACD & bcd  ; 
assign eid = ~EID;  //complement  
assign EIE =  ACA & ACB & ACC & ACD  ; 
assign eie = ~EIE;  //complement 
assign EIA =  ACA & bca  ; 
assign eia = ~EIA;  //complement 
assign EIB =  ACB & bcb  ; 
assign eib = ~EIB;  //complement 
assign EIC =  ACC & bcc  ; 
assign eic = ~EIC;  //complement 
assign acd = ~ACD;  //complement 
assign bcd = ~BCD;  //complement 
assign GJA = ~gja;  //complement 
assign GKA = ~gka;  //complement 
assign EJD =  ACH & bch  ; 
assign ejd = ~EJD;  //complement  
assign EJE =  ACE & ACF & ACG & ACH  ; 
assign eje = ~EJE;  //complement 
assign EJA =  ACE & bce  ; 
assign eja = ~EJA;  //complement 
assign EJB =  ACF & bcf  ; 
assign ejb = ~EJB;  //complement 
assign EJC =  ACG & bcg  ; 
assign ejc = ~EJC;  //complement 
assign ace = ~ACE;  //complement 
assign bce = ~BCE;  //complement 
assign JAJ =  GMD & HAE & QAE & HBE & HCA  |  ZZO & QAE & HBE & HCA  |  GED & HBE & HCA  |  GIA & HCA  |  GJA  ; 
assign jaj = ~JAJ;  //complement 
assign CJF =  ACE  ; 
assign cjf = ~CJF;  //complement 
assign CJG =  ACF & ACE  |  BCF  ; 
assign cjg = ~CJG;  //complement 
assign cje =  bce & bcf & bcg & bch  |  acf & bcg & bch  |  acg & bch  |  ach  ; 
assign CJE = ~cje;  //complement 
assign acf = ~ACF;  //complement 
assign bcf = ~BCF;  //complement 
assign kja = ~KJA;  //complement 
assign kje = ~KJE;  //complement 
assign CJH =  ACE & ACF & ACG  |  BCF & ACG  |  BCG  ; 
assign cjh = ~CJH;  //complement 
assign cjd =  bce & bcf & bcg  |  acf & bcg  |  acg  ; 
assign CJD = ~cjd;  //complement 
assign acg = ~ACG;  //complement 
assign bcg = ~BCG;  //complement 
assign kjc = ~KJC;  //complement 
assign kjg = ~KJG;  //complement 
assign cjb =  bce  ; 
assign CJB = ~cjb;  //complement 
assign cjc =  bcf & bce  |  acf  ; 
assign CJC = ~cjc;  //complement 
assign ach = ~ACH;  //complement 
assign bch = ~BCH;  //complement 
assign fga = ~FGA;  //complement 
assign fgb = ~FGB;  //complement 
assign fgc = ~FGC;  //complement 
assign fha = ~FHA;  //complement 
assign fhb = ~FHB;  //complement 
assign MAG =  kga & kgb & kgc & kgd  ; 
assign mag = ~MAG;  //complement  
assign MBG =  kge & kgf & kgg & kgh  ; 
assign mbg = ~MBG;  //complement 
assign NBH = ~nbh;  //complement 
assign MAH =  kha & khb & khc & khd  ; 
assign mah = ~MAH;  //complement  
assign MBH =  khe & khf & khg & khh  ; 
assign mbh = ~MBH;  //complement 
assign MDB =  KBE & KBF & KBG & KBH  ; 
assign mdb = ~MDB;  //complement  
assign MCG =  KGA & KGB & KGC & KGD  ; 
assign mcg = ~MCG;  //complement  
assign MDG =  KGE & KGF & KGG & KGH  ; 
assign mdg = ~MDG;  //complement 
assign kgb = ~KGB;  //complement 
assign kgf = ~KGF;  //complement 
assign sga =  kgc & KGB  |  KGD  ; 
assign SGA = ~sga;  //complement 
assign sgb =  KGC & kgb  |  kgd  ; 
assign SGB = ~sgb;  //complement 
assign fgd = ~FGD;  //complement 
assign kgh = ~KGH;  //complement 
assign kgd = ~KGD;  //complement 
assign sgc =  kgg & KGF  |  KGH  ; 
assign SGC = ~sgc;  //complement 
assign sgd =  KGG & kgf  |  kgh  ; 
assign SGD = ~sgd;  //complement 
assign NAG = ~nag;  //complement 
assign NBG = ~nbg;  //complement 
assign uga = ~UGA;  //complement 
assign ugb = ~UGB;  //complement 
assign pca =  naf & nbf  |  nag & nbg  |  nah & nbh  ; 
assign PCA = ~pca;  //complement 
assign pab =  nae & nbe  |  naf & nbf  |  nag & nbg  |  nah & nbh  ; 
assign PAB = ~pab;  //complement 
assign peb =  nae & nbe  |  naf & nbf  |  nag & nbg  |  nah & nbh  ; 
assign PEB = ~peb; //complement 
assign gmd = ~GMD;  //complement 
assign khb = ~KHB;  //complement 
assign pcc =  nah & nbh  |  NAG  |  NBG  ; 
assign PCC = ~pcc;  //complement 
assign pgc =  nah & nbh  |  NAG  |  NBG  ; 
assign PGC = ~pgc; //complement 
assign pcb =  NAF  |  NBF  |  nag & nbg  |  nah & nbh  ; 
assign PCB = ~pcb;  //complement 
assign pgb =  NAF  |  NBF  |  nag & nbg  |  nah & nbh  ; 
assign PGB = ~pgb; //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign shd =  KHG & khf  |  khh  ; 
assign SHD = ~shd;  //complement 
assign shc =  khg & KHF  |  KHH  ; 
assign SHC = ~shc;  //complement 
assign NAH = ~nah;  //complement 
assign uha = ~UHA;  //complement 
assign uhb = ~UHB;  //complement 
assign sha =  khc & KHB  |  KHD  ; 
assign SHA = ~sha;  //complement 
assign shb =  KHC & khb  |  khd  ; 
assign SHB = ~shb;  //complement 
assign khf = ~KHF;  //complement 
assign MCH =  KHA & KHB & KHC & KHD  ; 
assign mch = ~MCH;  //complement  
assign MDH =  KHE & KHF & KHG & KHH  ; 
assign mdh = ~MDH;  //complement 
assign fhc = ~FHC;  //complement 
assign fhd = ~FHD;  //complement 
assign khd = ~KHD;  //complement 
assign khh = ~KHH;  //complement 
assign kge = ~KGE;  //complement 
assign kga = ~KGA;  //complement 
assign cgb =  bbi  ; 
assign CGB = ~cgb;  //complement 
assign cgc =  bbj & bbi  |  abj  ; 
assign CGC = ~cgc;  //complement 
assign abi = ~ABI;  //complement 
assign bbi = ~BBI;  //complement 
assign kgc = ~KGC;  //complement 
assign kgg = ~KGG;  //complement 
assign CGF =  ABI  ; 
assign cgf = ~CGF;  //complement 
assign CGG =  ABJ & ABI  |  BBJ  ; 
assign cgg = ~CGG;  //complement 
assign cgd =  bbi & bbj & bbk  |  abj & bbk  |  abk  ; 
assign CGD = ~cgd;  //complement 
assign abj = ~ABJ;  //complement 
assign bbj = ~BBJ;  //complement 
assign JAG =  GIC & HCD & QAF & HAD & HBB  |  GMA & QAF & HAD & HBB  |  ZZO & HAD & HBB  |  GEC & HBB  |  GGA  ; 
assign jag = ~JAG;  //complement 
assign CGH =  ABI & ABJ & ABK  |  BBJ & ABK  |  BBK  ; 
assign cgh = ~CGH;  //complement 
assign cge =  bbi & bbj & bbk & bbl  |  abj & bbk & bbl  |  abk & bbl  |  abl  ; 
assign CGE = ~cge;  //complement 
assign abk = ~ABK;  //complement 
assign bbk = ~BBK;  //complement 
assign GHA = ~gha;  //complement 
assign EGD =  ABL & bbl  ; 
assign egd = ~EGD;  //complement  
assign EGE =  ABI & ABJ & ABK & ABL  ; 
assign ege = ~EGE;  //complement 
assign EGA =  ABI & bbi  ; 
assign ega = ~EGA;  //complement 
assign EGB =  ABJ & bbj  ; 
assign egb = ~EGB;  //complement 
assign EGC =  ABK & bbk  ; 
assign egc = ~EGC;  //complement 
assign abl = ~ABL;  //complement 
assign bbl = ~BBL;  //complement 
assign HCD = ~hcd;  //complement 
assign HCE = ~hce;  //complement 
assign EHD =  ABP & bbg  ; 
assign ehd = ~EHD;  //complement  
assign EHE =  ABM & ABN & ABO & ABP  ; 
assign ehe = ~EHE;  //complement 
assign EHA =  ABM & bbm  ; 
assign eha = ~EHA;  //complement 
assign EHB =  ABN & bbn  ; 
assign ehb = ~EHB;  //complement 
assign EHC =  ABO & bbo  ; 
assign ehc = ~EHC;  //complement 
assign abm = ~ABM;  //complement 
assign bbm = ~BBM;  //complement 
assign JAH =  GIB & HCE & QAE & HAE & HBC  |  GMD & QAE & HAE & HBC  |  ZZO & HAE & HBC  |  GED & HBC  |  GHA  ; 
assign jah = ~JAH;  //complement 
assign CHF =  ABM  ; 
assign chf = ~CHF;  //complement 
assign CHG =  ABN & ABM  |  BBN  ; 
assign chg = ~CHG;  //complement 
assign che =  bbm & bbn & bbo & bbp  |  abn & bbo & bbp  |  abo & bbp  |  abp  ; 
assign CHE = ~che;  //complement 
assign abn = ~ABN;  //complement 
assign bbn = ~BBN;  //complement 
assign kha = ~KHA;  //complement 
assign khe = ~KHE;  //complement 
assign CHH =  ABM & ABN & ABO  |  BBN & ABO  |  BBO  ; 
assign chh = ~CHH;  //complement 
assign chd =  bbm & bbn & bbo  |  abn & bbo  |  abo  ; 
assign CHD = ~chd;  //complement 
assign abo = ~ABO;  //complement 
assign bbo = ~BBO;  //complement 
assign khc = ~KHC;  //complement 
assign khg = ~KHG;  //complement 
assign chb =  bbm  ; 
assign CHB = ~chb;  //complement 
assign chc =  bbn & bbm  |  abn  ; 
assign CHC = ~chc;  //complement 
assign abp = ~ABP;  //complement 
assign bbp = ~BBP;  //complement 
assign MAE =  kea & keb & kec & ked  ; 
assign mae = ~MAE;  //complement  
assign MBE =  kee & kef & keg & keh  ; 
assign mbe = ~MBE;  //complement 
assign MAF =  kfa & kfb & kfc & kfd  ; 
assign maf = ~MAF;  //complement  
assign MBF =  kfe & kff & kfg & kfh  ; 
assign mbf = ~MBF;  //complement 
assign MCE =  KEA & KEB & KEC & KED  ; 
assign mce = ~MCE;  //complement  
assign MDE =  KEE & KEF & KEG & KEH  ; 
assign mde = ~MDE;  //complement 
assign fea = ~FEA;  //complement 
assign feb = ~FEB;  //complement 
assign keb = ~KEB;  //complement 
assign kef = ~KEF;  //complement 
assign sea =  kec & KEB  |  KED  ; 
assign SEA = ~sea;  //complement 
assign seb =  KEC & keb  |  ked  ; 
assign SEB = ~seb;  //complement 
assign fec = ~FEC;  //complement 
assign fed = ~FED;  //complement 
assign ked = ~KED;  //complement 
assign keh = ~KEH;  //complement 
assign sed =  KEG & kef  |  keh  ; 
assign SED = ~sed;  //complement 
assign sec =  keg & KEF  |  KEH  ; 
assign SEC = ~sec;  //complement 
assign ffa = ~FFA;  //complement 
assign ffb = ~FFB;  //complement 
assign NAE = ~nae;  //complement 
assign NBE = ~nbe;  //complement 
assign uea = ~UEA;  //complement 
assign ueb = ~UEB;  //complement 
assign pbd =  NAD  |  NBD  ; 
assign PBD = ~pbd;  //complement 
assign gmc = ~GMC;  //complement 
assign oia = ~OIA;  //complement 
assign gea = ~GEA;  //complement 
assign sfc =  kfg & KFF  |  KFH  ; 
assign SFC = ~sfc;  //complement 
assign sfd =  KFG & kff  |  kfh  ; 
assign SFD = ~sfd;  //complement 
assign NAF = ~naf;  //complement 
assign NBF = ~nbf;  //complement 
assign ufa = ~UFA;  //complement 
assign ufb = ~UFB;  //complement 
assign sfa =  kfc & KFB  |  KFD  ; 
assign SFA = ~sfa;  //complement 
assign sfb =  KFC & kfb  |  kfd  ; 
assign SFB = ~sfb;  //complement 
assign kfb = ~KFB;  //complement 
assign kff = ~KFF;  //complement 
assign MCF =  KFA & KFB & KFC & KFD  ; 
assign mcf = ~MCF;  //complement  
assign MDF =  KFE & KFF & KFG & KFH  ; 
assign mdf = ~MDF;  //complement 
assign ffc = ~FFC;  //complement 
assign ffd = ~FFD;  //complement 
assign kfd = ~KFD;  //complement 
assign kfh = ~KFH;  //complement 
assign kea = ~KEA;  //complement 
assign kee = ~KEE;  //complement 
assign ceb =  bba  ; 
assign CEB = ~ceb;  //complement 
assign cec =  bbb & bba  |  abb  ; 
assign CEC = ~cec;  //complement 
assign aba = ~ABA;  //complement 
assign bba = ~BBA;  //complement 
assign kec = ~KEC;  //complement 
assign keg = ~KEG;  //complement 
assign CEF =  ABA  ; 
assign cef = ~CEF;  //complement 
assign CEG =  ABB & ABA  |  BBB  ; 
assign ceg = ~CEG;  //complement 
assign ced =  bba & bbb & bbc  |  abb & bbc  |  abc  ; 
assign CED = ~ced;  //complement 
assign abb = ~ABB;  //complement 
assign bbb = ~BBB;  //complement 
assign JAE =  GIC & HCD & HAD & QAD  |  GMC & HAD & QAD  |  GEA & QAD  ; 
assign jae = ~JAE;  //complement 
assign CEH =  ABA & ABB & ABC  |  BBB & ABC  |  BBC  ; 
assign ceh = ~CEH;  //complement 
assign cee =  bba & bbb & bbc & bbd  |  abb & bbc & bbd  |  abc & bbd  |  abd  ; 
assign CEE = ~cee;  //complement 
assign abc = ~ABC;  //complement 
assign bbc = ~BBC;  //complement 
assign GFA = ~gfa;  //complement 
assign GGA = ~gga;  //complement 
assign EED =  ABD & bbd  ; 
assign eed = ~EED;  //complement  
assign EEE =  ABA & ABB & ABC & ABD  ; 
assign eee = ~EEE;  //complement 
assign EEA =  ABA & bba  ; 
assign eea = ~EEA;  //complement 
assign EEB =  ABB & bbb  ; 
assign eeb = ~EEB;  //complement 
assign EEC =  ABC & bbc  ; 
assign eec = ~EEC;  //complement 
assign abd = ~ABD;  //complement 
assign bbd = ~BBD;  //complement 
assign GLA = ~gla;  //complement 
assign EFD =  ABH & bbh  ; 
assign efd = ~EFD;  //complement  
assign EFE =  ABE & ABF & ABG & ABH  ; 
assign efe = ~EFE;  //complement 
assign EFA =  ABE & bbe  ; 
assign efa = ~EFA;  //complement 
assign EFB =  ABF & bbf  ; 
assign efb = ~EFB;  //complement 
assign EFC =  ABG & bbg  ; 
assign efc = ~EFC;  //complement 
assign abe = ~ABE;  //complement 
assign bbe = ~BBE;  //complement 
assign JAF =  GIB & HCE & QAC & HAE & HBA  |  GMB & QAC & HAE & HBA  |  ZZO & HAE & HBA  |  GED & HBA  |  GFA  ; 
assign jaf = ~JAF;  //complement 
assign CFF =  ABE  ; 
assign cff = ~CFF;  //complement 
assign CFG =  ABF & ABE  |  BBF  ; 
assign cfg = ~CFG;  //complement 
assign cfe =  bbe & bbf & bbg & bbh  |  abf & bbg & bbh  |  abg & bbh  |  abh  ; 
assign CFE = ~cfe;  //complement 
assign abf = ~ABF;  //complement 
assign bbf = ~BBF;  //complement 
assign kfa = ~KFA;  //complement 
assign kfe = ~KFE;  //complement 
assign CFH =  ABE & ABF & ABG  |  BBF & ABG  |  BBG  ; 
assign cfh = ~CFH;  //complement 
assign sja =  kjc & KJB  |  KJD  ; 
assign SJA = ~sja;  //complement 
assign abg = ~ABG;  //complement 
assign bbg = ~BBG;  //complement 
assign kfc = ~KFC;  //complement 
assign kfg = ~KFG;  //complement 
assign cfd =  bbe & bbf & bbg  |  abf & bbg  |  abg  ; 
assign CFD = ~cfd;  //complement 
assign cfb =  bbe  ; 
assign CFB = ~cfb;  //complement 
assign cfc =  bbf & bbe  |  abf  ; 
assign CFC = ~cfc;  //complement 
assign abh = ~ABH;  //complement 
assign bbh = ~BBH;  //complement 
assign MAC =  kca & kcb & kcc & kcd  ; 
assign mac = ~MAC;  //complement  
assign MBC =  kce & kcf & kcg & kch  ; 
assign mbc = ~MBC;  //complement 
assign MAD =  kda & kdb & kdc & kdd  ; 
assign mad = ~MAD;  //complement  
assign MBD =  kde & kdf & kdg & kdh  ; 
assign mbd = ~MBD;  //complement 
assign MCC =  KCA & KCB & KCC & KCD  ; 
assign mcc = ~MCC;  //complement  
assign MDC =  KCE & KCF & KCG & KCH  ; 
assign mdc = ~MDC;  //complement 
assign fca = ~FCA;  //complement 
assign fcb = ~FCB;  //complement 
assign kcb = ~KCB;  //complement 
assign kcf = ~KCF;  //complement 
assign sca =  kcc & KCB  |  KCD  ; 
assign SCA = ~sca;  //complement 
assign scb =  KCC & kcb  |  kcd  ; 
assign SCB = ~scb;  //complement 
assign fcc = ~FCC;  //complement 
assign fcd = ~FCD;  //complement 
assign kcd = ~KCD;  //complement 
assign kch = ~KCH;  //complement 
assign scc =  kcg & KCF  |  KCH  ; 
assign SCC = ~scc;  //complement 
assign scd =  KCG & kcf  |  kch  ; 
assign SCD = ~scd;  //complement 
assign fda = ~FDA;  //complement 
assign fdb = ~FDB;  //complement 
assign NAC = ~nac;  //complement 
assign NBC = ~nbc;  //complement 
assign uca = ~UCA;  //complement 
assign ucb = ~UCB;  //complement 
assign pba =  nab & nbb  |  nac & nbc  |  nad & nbd  ; 
assign PBA = ~pba;  //complement 
assign paa =  naa & nba  |  nab & nbb  |  nac & nbc  |  nad & nbd  ; 
assign PAA = ~paa;  //complement 
assign gma = ~GMA;  //complement 
assign pbc =  NAC  |  NBC  |  nad & nbd  ; 
assign PBC = ~pbc;  //complement 
assign pfc =  NAC  |  NBC  |  nad & nbd  ; 
assign PFC = ~pfc; //complement 
assign pbb =  NAB  |  NBB  |  nac & nbc  |  nad & nbd  ; 
assign PBB = ~pbb;  //complement 
assign pfb =  NAB  |  NBB  |  nac & nbc  |  nad & nbd  ; 
assign PFB = ~pfb; //complement 
assign sdc =  kdg & KDF  |  KDH  ; 
assign SDC = ~sdc;  //complement 
assign sdd =  KDG & kdf  |  kdh  ; 
assign SDD = ~sdd;  //complement 
assign NAD = ~nad;  //complement 
assign NBD = ~nbd;  //complement 
assign uda = ~UDA;  //complement 
assign udb = ~UDB;  //complement 
assign sda =  kdc & KDB  |  KDD  ; 
assign SDA = ~sda;  //complement 
assign sdb =  KDC & kdb  |  kdd  ; 
assign SDB = ~sdb;  //complement 
assign kdb = ~KDB;  //complement 
assign kdf = ~KDF;  //complement 
assign MCD =  KDA & KDB & KDC & KDD  ; 
assign mcd = ~MCD;  //complement  
assign MDD =  KDE & KDF & KDG & KDH  ; 
assign mdd = ~MDD;  //complement 
assign fdc = ~FDC;  //complement 
assign fdd = ~FDD;  //complement 
assign kdd = ~KDD;  //complement 
assign kdh = ~KDH;  //complement 
assign kca = ~KCA;  //complement 
assign kce = ~KCE;  //complement 
assign GDA = ~gda;  //complement 
assign ccb =  bai  ; 
assign CCB = ~ccb;  //complement 
assign ccc =  baj & bai  |  aai  ; 
assign CCC = ~ccc;  //complement 
assign aai = ~AAI;  //complement 
assign bai = ~BAI;  //complement 
assign kcc = ~KCC;  //complement 
assign kcg = ~KCG;  //complement 
assign CCF =  AAI  ; 
assign ccf = ~CCF;  //complement 
assign CCG =  AAJ & AAI  |  BAJ  ; 
assign ccg = ~CCG;  //complement 
assign ccd =  bai & baj & bak  |  aaj & bak  |  aak  ; 
assign CCD = ~ccd;  //complement 
assign aaj = ~AAJ;  //complement 
assign baj = ~BAJ;  //complement 
assign JAC =  GEA & HBD & HCD & HAB & QAD  |  GID & HCD & HAB & QAD  |  GMC & HAB & QAD  |  GCA & QAD  ; 
assign jac = ~JAC;  //complement 
assign CCH =  AAI & AAJ & AAK  |  BAJ & AAK  |  BAK  ; 
assign cch = ~CCH;  //complement 
assign cce =  bai & baj & bak & bal  |  aaj & bak & bal  |  aak & bal  |  aal  ; 
assign CCE = ~cce;  //complement 
assign aak = ~AAK;  //complement 
assign bak = ~BAK;  //complement 
assign ECD =  AAL & bal  ; 
assign ecd = ~ECD;  //complement  
assign ECE =  AAI & AAJ & AAK & AAL  ; 
assign ece = ~ECE;  //complement 
assign ECA =  AAI & bai  ; 
assign eca = ~ECA;  //complement 
assign ECB =  AAJ & baj  ; 
assign ecb = ~ECB;  //complement 
assign ECC =  AAK & bak  ; 
assign ecc = ~ECC;  //complement 
assign aal = ~AAL;  //complement 
assign bal = ~BAL;  //complement 
assign bao = ~BAO;  //complement 
assign EDE =  AAM & AAN & AAO & AAP  ; 
assign ede = ~EDE;  //complement  
assign EDD =  AAP & bap  ; 
assign edd = ~EDD;  //complement 
assign EDA =  AAM & bam  ; 
assign eda = ~EDA;  //complement 
assign EDB =  AAN & ban  ; 
assign edb = ~EDB;  //complement 
assign EDC =  AAO & bao  ; 
assign edc = ~EDC;  //complement 
assign aam = ~AAM;  //complement 
assign bam = ~BAM;  //complement 
assign JAD =  GEB & HBE & HCE & HAC & QAC  |  GIA & HCE & HAC & QAC  |  GMB & HAC & QAC  |  GDA & QAC  ; 
assign jad = ~JAD;  //complement 
assign CDF =  AAM  ; 
assign cdf = ~CDF;  //complement 
assign CDG =  AAN & AAM  |  BAN  ; 
assign cdg = ~CDG;  //complement 
assign cde =  bam & ban & bao & bap  |  aan & bao & bap  |  aao & bap  |  aap  ; 
assign CDE = ~cde;  //complement 
assign aan = ~AAN;  //complement 
assign ban = ~BAN;  //complement 
assign kda = ~KDA;  //complement 
assign kde = ~KDE;  //complement 
assign CDH =  AAM & AAN & AAO  |  BAN & AAO  |  BAO  ; 
assign cdh = ~CDH;  //complement 
assign cdd =  bam & ban & bao  |  aan & bao  |  aao  ; 
assign CDD = ~cdd;  //complement 
assign aao = ~AAO;  //complement 
assign kdc = ~KDC;  //complement 
assign kdg = ~KDG;  //complement 
assign cdb =  bam  ; 
assign CDB = ~cdb;  //complement 
assign cdc =  ban & bam  |  aan  ; 
assign CDC = ~cdc;  //complement 
assign aap = ~AAP;  //complement 
assign bap = ~BAP;  //complement 
assign MAA =  kaa & kab & kac & kad  ; 
assign maa = ~MAA;  //complement  
assign MBA =  kae & kaf & kag & kah  ; 
assign mba = ~MBA;  //complement 
assign MAB =  kba & kbb & kbc & kbd  ; 
assign mab = ~MAB;  //complement  
assign MBB =  kbe & kbf & kbg & kbh  ; 
assign mbb = ~MBB;  //complement 
assign MCA =  KAA & KAB & KAC & KAD  ; 
assign mca = ~MCA;  //complement  
assign MDA =  KAE & KAF & KAG & KAH  ; 
assign mda = ~MDA;  //complement 
assign faa = ~FAA;  //complement 
assign fab = ~FAB;  //complement 
assign kab = ~KAB;  //complement 
assign kaf = ~KAF;  //complement 
assign saa =  kac & KAB  |  KAD  ; 
assign SAA = ~saa;  //complement 
assign sab =  KAC & kab  |  kad  ; 
assign SAB = ~sab;  //complement 
assign fac = ~FAC;  //complement 
assign fad = ~FAD;  //complement 
assign kad = ~KAD;  //complement 
assign kah = ~KAH;  //complement 
assign sac =  kag & KAF  |  KAH  ; 
assign SAC = ~sac;  //complement 
assign sad =  KAG & kaf  |  kah  ; 
assign SAD = ~sad;  //complement 
assign fba = ~FBA;  //complement 
assign fbb = ~FBB;  //complement 
assign NAA = ~naa;  //complement 
assign uaa = ~UAA;  //complement 
assign uab = ~UAB;  //complement 
assign gmb = ~GMB;  //complement 
assign kbb = ~KBB;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign sbc =  kbg & KBF  |  KBH  ; 
assign SBC = ~sbc;  //complement 
assign sbd =  KBG & kbf  |  kbh  ; 
assign SBD = ~sbd;  //complement 
assign NBA = ~nba;  //complement 
assign NAB = ~nab;  //complement 
assign NBB = ~nbb;  //complement 
assign uba = ~UBA;  //complement 
assign ubb = ~UBB;  //complement 
assign sba =  kbc & KBB  |  KBD  ; 
assign SBA = ~sba;  //complement 
assign sbb =  KBC & kbb  |  kbd  ; 
assign SBB = ~sbb;  //complement 
assign kbf = ~KBF;  //complement 
assign MCB =  KBA & KBB & KBC & KBD  ; 
assign mcb = ~MCB;  //complement  
assign fbc = ~FBC;  //complement 
assign fbd = ~FBD;  //complement 
assign kbd = ~KBD;  //complement 
assign kbh = ~KBH;  //complement 
assign kaa = ~KAA;  //complement 
assign kae = ~KAE;  //complement 
assign kba = ~KBA;  //complement 
assign aaa = ~AAA;  //complement 
assign AAR = ~aar;  //complement 
assign cab =  baa  ; 
assign CAB = ~cab;  //complement 
assign cac =  bab & baa  |  aab  ; 
assign CAC = ~cac;  //complement 
assign aaq = ~AAQ;  //complement 
assign BAA = ~baa;  //complement 
assign kac = ~KAC;  //complement 
assign kag = ~KAG;  //complement 
assign CAF =  AAA  ; 
assign caf = ~CAF;  //complement 
assign CAG =  AAB & AAA  |  BAB  ; 
assign cag = ~CAG;  //complement 
assign fid = ~FID;  //complement 
assign aab = ~AAB;  //complement 
assign bab = ~BAB;  //complement 
assign JAA =  GEA & HBD & HCD & QAD  |  GID & HCD & QAD  |  GMC & QAD  ; 
assign jaa = ~JAA;  //complement 
assign CAH =  AAA & AAB & AAC  |  BAB & AAC  |  BAC  ; 
assign cah = ~CAH;  //complement 
assign cad =  baa & bab & bac  |  aab & bac  |  aac  ; 
assign CAD = ~cad;  //complement 
assign aac = ~AAC;  //complement 
assign bac = ~BAC;  //complement 
assign GBA = ~gba;  //complement 
assign EAD =  AAD & bad  ; 
assign ead = ~EAD;  //complement  
assign EAE =  AAB & AAC & AAD  ; 
assign eae = ~EAE;  //complement 
assign EAA =  AAQ  ; 
assign eaa = ~EAA;  //complement 
assign EAB =  AAB & bab  ; 
assign eab = ~EAB;  //complement 
assign EAC =  AAC & bac  ; 
assign eac = ~EAC;  //complement 
assign aad = ~AAD;  //complement 
assign bad = ~BAD;  //complement 
assign HCA = ~hca;  //complement 
assign HCB = ~hcb;  //complement 
assign EBD =  AAH & bah  ; 
assign ebd = ~EBD;  //complement  
assign EBE =  AAE & AAF & AAG & AAH  ; 
assign ebe = ~EBE;  //complement 
assign EBA =  AAE & bae  ; 
assign eba = ~EBA;  //complement 
assign EBB =  AAF & baf  ; 
assign ebb = ~EBB;  //complement 
assign EBC =  AAG & bag  ; 
assign ebc = ~EBC;  //complement 
assign aae = ~AAE;  //complement 
assign bae = ~BAE;  //complement 
assign JAB =  GEB & HBE & HCE & HAA & QAC  |  GIA & HCE & HAA & QAC  |  GMB & HAA & QAC  |  GBA & QAC  ; 
assign jab = ~JAB;  //complement 
assign CBF =  AAE  ; 
assign cbf = ~CBF;  //complement 
assign CBG =  AAF & AAE  |  BAF  ; 
assign cbg = ~CBG;  //complement 
assign cbe =  bae & baf & bag & bah  |  aaf & bag & bah  |  aag & bah  |  aah  ; 
assign CBE = ~cbe;  //complement 
assign aaf = ~AAF;  //complement 
assign baf = ~BAF;  //complement 
assign kbe = ~KBE;  //complement 
assign CBH =  AAE & AAF & AAG  |  BAF & AAG  |  BAG  ; 
assign cbh = ~CBH;  //complement 
assign cbd =  bae & baf & bag  |  aaf & bag  |  aag  ; 
assign CBD = ~cbd;  //complement 
assign aag = ~AAG;  //complement 
assign bag = ~BAG;  //complement 
assign kbc = ~KBC;  //complement 
assign kbg = ~KBG;  //complement 
assign cae =  baa & bab & bac & bad  |  aab & bac & bad  |  aac & bad  |  aad  ; 
assign CAE = ~cae;  //complement 
assign cbb =  bae  ; 
assign CBB = ~cbb;  //complement 
assign cbc =  baf & bae  |  aaf  ; 
assign CBC = ~cbc;  //complement 
assign aah = ~AAH;  //complement 
assign bah = ~BAH;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iar = ~IAR; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibm = ~IBM; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iff = ~IFF; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
always@(posedge IZZ )
   begin 
 QDA <= JAM & QAH ; 
 QDB <= JAM & qah ; 
 GID <=  CEE & EFE & EGE & EHE  |  CFE & EGE & EHE  |  CGE & EHE  |  CHE  ; 
 oha <= qda ; 
 qga <= qca ; 
 gca <=  cae & cbe  |  ebe & cbe  ; 
 OHB <= qga & QDB ; 
 OCA <= FIA & qbb |  fia & QBB ; 
 OCB <= FIB & qbb |  fib & QBB ; 
 OCC <= FIC & qbb |  fic & QBB ; 
 OBI <= FGA & qbb |  fga & QBB ; 
 OBJ <= FGB & qbb |  fgb & QBB ; 
 OCD <= FID & qbb |  fid & QBB ; 
 qbe <= jbc ; 
 qbf <= jbc ; 
 qbg <= jbc ; 
 qbh <= jbc ; 
 ode <=  ZZO & PEB & PEC  |  ZZO & PEB & PEC  |  pba & PEB & PEC  |  pca & peb & PEC  |  pda & pec  ; 
 OBK <= FGC & qbb |  fgc & QBB ; 
 OBL <= FGD & qbb |  fgd & QBB ; 
 OCI <= FKA & qbb |  fka & QBB ; 
 qba <= jbc ; 
 qbb <= jbc ; 
 qbc <= jbc ; 
 qbd <= jbc ; 
 OFA <=  REA & PCA  |  RFA & PCB  |  RGA & PCC  |  RHA & PCD  ; 
 OGA <=  RIA & PDA  |  RJA & PDB  |  RKA & PDC  |  RLA & PDD  ; 
 OCJ <= FKB & qbb |  fkb & QBB ; 
 OCK <= FKC & qbb |  fkc & QBB ; 
 OCL <= FKD & qbb |  fkd & QBB ; 
 haa <=  eae  ; 
 hab <=  eae  |  ebe  ; 
 OEA <=  RAA & PBA  |  RBA & PBB  |  RCA & PBC  |  RDA & PBD  ; 
 ODC <=  ZZO & PEB & PEC  |  ZZO & PEB & PEC  |  PFB & PEB & PEC  |  PGB & peb & PEC  |  PHB & pec  ; 
 OCM <= FLA & qbc |  fla & QBC ; 
 OCN <= FLB & qbc |  flb & QBC ; 
 OCO <= FLC & qbc |  flc & QBC ; 
 OBM <= FHA & qbc |  fha & QBC ; 
 OBN <= FHB & qbc |  fhb & QBC ; 
 OCP <= FLD & qbc |  fld & QBC ; 
 OBO <= FHC & qbc |  fhc & QBC ; 
 OBP <= FHD & qbc |  fhd & QBC ; 
 OCE <= FJA & qbc |  fja & QBC ; 
 OCF <= FJB & qbc |  fjb & QBC ; 
 OCG <= FJC & qbc |  fjc & QBC ; 
 OCH <= FJD & qbc |  fjd & QBC ; 
 QAB <= IJA ; 
 QCA <= QAB & qaa ; 
 QFA <= QAB & QAB ; 
 QAA <= IJA & IJB ; 
 GIC <=  CEE & EFE & EGE & EHE  |  CFE & EGE & EHE  |  CGE & EHE  |  CHE  ; 
 QAG <= QAA ; 
 QAH <= QAA ; 
 GEC <=  CAE & EBE & ECE & EDE  |  CBE & ECE & EDE  |  CCE & EDE  |  CDE  ; 
 OAI <= FCA & qba |  fca & QBA ; 
 OAJ <= FCB & qba |  fcb & QBA ; 
 OAK <= FCC & qba |  fcc & QBA ; 
 OAA <= FAA & qba |  faa & QBA ; 
 OAB <= FAB & qba |  fab & QBA ; 
 OAL <= FCD & qba |  fcd & QBA ; 
 OAC <= FAC & qba |  fac & QBA ; 
 OAD <= FAD & qba |  fad & QBA ; 
 OBA <= FEA & qba |  fea & QBA ; 
 hba <=  eee  ; 
 hbb <=  eee  |  efe  ; 
 OFB <=  REB & PCA  |  RFB & PCB  |  RGB & PCC  |  RHB & PCD  ; 
 OGB <=  RIB & PDA  |  RJB & PDB  |  RKB & PDC  |  RLB & PDD  ; 
 OBB <= FEB & qba |  feb & QBA ; 
 OBC <= FEC & qba |  fec & QBA ; 
 OBD <= FED & qba |  fed & QBA ; 
 hac <=  eae  |  ebe  |  ece  ; 
 OEB <=  RAB & PBA  |  RBB & PBB  |  RCB & PBC  |  RDB & PBD  ; 
 ODD <=  ZZO & PEB & PEC  |  ZZO & PEB & PEC  |  PFC & PEB & PEC  |  PGC & peb & PEC  |  PHC & pec  ; 
 OBE <= FFA & qbd |  ffa & QBD ; 
 OBF <= FFB & qbd |  ffb & QBD ; 
 OBG <= FFC & qbd |  ffc & QBD ; 
 QFB <= QFA ; 
 ojb <= qfb ; 
 oja <= qec ; 
 qea <= ijb ; 
 qeb <= qea ; 
 qec <= qeb ; 
 OAE <= FBA & qbd |  fba & QBD ; 
 OAF <= FBB & qbd |  fbb & QBD ; 
 OBH <= FFD & qbd |  ffd & QBD ; 
 OAG <= FBC & qbd |  fbc & QBD ; 
 OAH <= FBD & qbd |  fbd & QBD ; 
 OAM <= FDA & qbd |  fda & QBD ; 
 OAN <= FDB & qbd |  fdb & QBD ; 
 OAO <= FDC & qbd |  fdc & QBD ; 
 OAP <= FDD & qbd |  fdd & QBD ; 
 FKA <=  KKA & jak  |  KKE & JAK  ; 
 FKB <=  KKB & jak  |  KKF & JAK  ; 
 KKB <=  ckb & EKB  |  CKB & ekb  ; 
 KKF <=  ckf & EKB  |  CKF & ekb  ; 
 FKC <=  KKC & jak  |  KKG & JAK  ; 
 FKD <=  KKD & jak  |  KKH & JAK  ; 
 KKD <=  ckd & EKD  |  CKD & ekd  ; 
 KKH <=  ckh & EKD  |  CKH & ekd  ; 
 FLA <=  KLA & jal  |  KLE & JAL  ; 
 FLB <=  KLB & jal  |  KLF & JAL  ; 
 nak <=  mak & jak  |  mbk & JAK  |  JBB  ; 
 nbk <=  mck & jak  |  mdk & JAK  |  jbb  ; 
 UKA <=  SKA & jak  |  SKC & JAK  ; 
 UKB <=  SKB & jak  |  SKD & JAK  ; 
 GIB <=  CEE & EFE & EGE & EHE  |  CFE & EGE & EHE  |  CGE & EHE  |  CHE  ; 
 GED <=  CAE & EBE & ECE & EDE  |  CBE & ECE & EDE  |  CCE & EDE  |  CDE  ; 
 nal <=  mal & jal  |  mbl & JAL  |  JBA  ; 
 nbl <=  mcl & jal  |  mdl & JAL  |  jba  ; 
 ULA <=  SLA & jal  |  SLC & JAL  ; 
 ULB <=  SLB & jal  |  SLD & JAL  ; 
 KLB <=  clb & ELB  |  CLB & elb  ; 
 KLF <=  clf & ELB  |  CLF & elb  ; 
 FLC <=  KLC & jal  |  KLG & JAL  ; 
 FLD <=  KLD & jal  |  KLH & JAL  ; 
 KLD <=  cld & ELD  |  CLD & eld  ; 
 KLH <=  clh & ELD  |  CLH & eld  ; 
 KKA <=  EKA  ; 
 KKE <=  eka  ; 
 ACI <=  IFI & IFI  |  ICI  ; 
 BCI <=  ICI & IFI  ; 
 KKC <=  ckc & EKC  |  CKC & ekc  ; 
 KKG <=  ckg & EKC  |  CKG & ekc  ; 
 ACJ <=  IFJ & IFJ  |  ICJ  ; 
 BCJ <=  ICJ & IFJ  ; 
 ACK <=  IFK & IFK  |  ICK  ; 
 BCK <=  ICK & IFK  ; 
 hbd <=  eee  |  efe  |  ege  |  ehe  ; 
 hbe <=  eee  |  efe  |  ege  |  ehe  ; 
 ACL <=  IFL & IFL  |  ICL  ; 
 BCL <=  ICL & IFL  ; 
 had <=  eae  |  ebe  |  ece  |  ede  ; 
 hae <=  eae  |  ebe  |  ece  |  ede  ; 
 ACM <=  IFM & IFM  |  ICM  ; 
 BCM <=  ICM & IFM  ; 
 ACN <=  IFN & IFN  |  ICN  ; 
 BCN <=  ICN & IFN  ; 
 KLA <=  ELA  ; 
 KLE <=  ela  ; 
 ACO <=  IFO & IFO  |  ICO  ; 
 BCO <=  ICO & IFO  ; 
 KLC <=  clc & ELC  |  CLC & elc  ; 
 KLG <=  clg & ELC  |  CLG & elc  ; 
 ACP <=  IFP & IFP  |  ICP  ; 
 BCP <=  ICP & IFP  ; 
 FIA <=  KIA & jai  |  KIE & JAI  ; 
 FIB <=  KIB & jai  |  KIF & JAI  ; 
 KIB <=  cib & EIB  |  CIB & eib  ; 
 KIF <=  cif & EIB  |  CIF & eib  ; 
 FIC <=  KIC & jai  |  KIG & JAI  ; 
 KID <=  cid & EID  |  CID & eid  ; 
 KIH <=  cih & EID  |  CIH & eid  ; 
 FJA <=  KJA & jaj  |  KJE & JAJ  ; 
 FJB <=  KJB & jaj  |  KJF & JAJ  ; 
 nai <=  mai & jai  |  mbi & JAI  |  JBB  ; 
 nbi <=  mci & jai  |  mdi & JAI  |  jbb  ; 
 UIA <=  SIA & jai  |  SIC & JAI  ; 
 UIB <=  SIB & jai  |  SID & JAI  ; 
 GIA <=  CEE & EFE & EGE & EHE  |  CFE & EGE & EHE  |  CGE & EHE  |  CHE  ; 
 KJB <=  cjb & EJB  |  CJB & ejb  ; 
 KJF <=  cjf & EJB  |  CJF & ejb  ; 
 GEB <=  CAE & EBE & ECE & EDE  |  CBE & ECE & EDE  |  CCE & EDE  |  CDE  ; 
 naj <=  maj & jaj  |  mbj & JAJ  |  JBA  ; 
 nbj <=  mcj & jaj  |  mdj & JAJ  |  jba  ; 
 UJA <=  SJA & jaj  |  SJC & JAJ  ; 
 UJB <=  SJB & jaj  |  SJD & JAJ  ; 
 FJC <=  KJC & jaj  |  KJG & JAJ  ; 
 FJD <=  KJD & jaj  |  KJH & JAJ  ; 
 KJD <=  cjd & EJD  |  CJD & ejd  ; 
 KJH <=  cjh & EJD  |  CJH & ejd  ; 
 KIA <=  EIA  ; 
 KIE <=  eia  ; 
 ACA <=  IFA & IFA  |  ICA  ; 
 BCA <=  ICA & IFA  ; 
 KIC <=  cic & EIC  |  CIC & eic  ; 
 KIG <=  cig & EIC  |  CIG & eic  ; 
 ACB <=  IFB & IFB  |  ICB  ; 
 BCB <=  ICB & IFB  ; 
 ACC <=  IFC & IFC  |  ICC  ; 
 BCC <=  ICC & IFC  ; 
 hbc <=  eee  |  efe  |  ege  ; 
 hcc <=  eie  |  eje  |  eke  ; 
 ACD <=  IFD & IFD  |  ICD  ; 
 BCD <=  ICD & IFD  ; 
 gja <=  cie & cie  ; 
 gka <=  cje & cie  |  cie & eje  ; 
 ACE <=  IFE & IFE  |  ICE  ; 
 BCE <=  ICE & IFE  ; 
 ACF <=  IFF & IFF  |  ICF  ; 
 BCF <=  ICF & IFF  ; 
 KJA <=  EJA  ; 
 KJE <=  eja  ; 
 ACG <=  IFG & IFG  |  ICG  ; 
 BCG <=  ICG & IFG  ; 
 KJC <=  cjc & EJC  |  CJC & ejc  ; 
 KJG <=  cjg & EJC  |  CJG & ejc  ; 
 ACH <=  IFH & IFH  |  ICH  ; 
 BCH <=  ICH & IFH  ; 
 FGA <=  KGA & jag  |  KGE & JAG  ; 
 FGB <=  KGB & jag  |  KGF & JAG  ; 
 FGC <=  KGC & jag  |  KGG & JAG  ; 
 FHA <=  KHA & jah  |  KHE & JAH  ; 
 FHB <=  KHB & jah  |  KHF & JAH  ; 
 nbh <=  mch & jah  |  mdh & JAH  |  jba  ; 
 KGB <=  cgb & EGB  |  CGB & egb  ; 
 KGF <=  cgf & EGB  |  CGF & egb  ; 
 FGD <=  KGD & jag  |  KGH & JAG  ; 
 KGH <=  cgh & EGD  |  CGH & egd  ; 
 KGD <=  cgd & EGD  |  CGD & egd  ; 
 nag <=  mag & jag  |  mbg & JAG  |  JBB  ; 
 nbg <=  mcg & jag  |  mdg & JAG  |  jbb  ; 
 UGA <=  SGA & jag  |  SGC & JAG  ; 
 UGB <=  SGB & jag  |  SGD & JAG  ; 
 GMD <=  CIE & EJE & EKE & ELE  |  CJE & EKE & ELE  |  CKE & ELE  |  CLE  ; 
 KHB <=  chb & EHB  |  CHB & ehb  ; 
 QAC <= aar & QAA ; 
 QAD <= aar & QAA ; 
 QAE <= aar & QAA ; 
 QAF <= aar & QAA ; 
 nah <=  mah & jah  |  mbh & JAH  |  JBA  ; 
 UHA <=  SHA & jah  |  SHC & JAH  ; 
 UHB <=  SHB & jah  |  SHD & JAH  ; 
 KHF <=  chf & EHB  |  CHF & ehb  ; 
 FHC <=  KHC & jah  |  KHG & JAH  ; 
 FHD <=  KHD & jah  |  KHH & JAH  ; 
 KHD <=  chd & EHD  |  CHD & ehd  ; 
 KHH <=  chh & EHD  |  CHH & ehd  ; 
 KGE <=  ega  ; 
 KGA <=  EGA  ; 
 ABI <=  IEI & IEI  |  IBI  ; 
 BBI <=  IBI & IEI  ; 
 KGC <=  cgc & EGC  |  CGC & egc  ; 
 KGG <=  cgg & EGC  |  CGG & egc  ; 
 ABJ <=  IEJ & IEJ  |  IBJ  ; 
 BBJ <=  IBJ & IEJ  ; 
 ABK <=  IEK & IEK  |  IBK  ; 
 BBK <=  IBK & IEK  ; 
 gha <=  ZZO & cee & cfe & cge  |  ZZI & cee & cfe & cge  |  efe & cfe & cge  |  ege & cge & cge  ; 
 ABL <=  IEL & IEL  |  IBL  ; 
 BBL <=  IBL & IEL  ; 
 hcd <=  eie  |  eje  |  eke  |  ele  ; 
 hce <=  eie  |  eje  |  eke  |  ele  ; 
 ABM <=  IEM & IEM  |  IBM  ; 
 BBM <=  IBM & IEM  ; 
 ABN <=  IEN & IEN  |  IBN  ; 
 BBN <=  IBN & IEN  ; 
 KHA <=  EHA  ; 
 KHE <=  eha  ; 
 ABO <=  IEO & IEO  |  IBO  ; 
 BBO <=  IBO & IEO  ; 
 KHC <=  chc & EHC  |  CHC & ehc  ; 
 KHG <=  chg & EHC  |  CHG & ehc  ; 
 ABP <=  IEP & IEP  |  IBP  ; 
 BBP <=  IBP & IEP  ; 
 FEA <=  KEA & jae  |  KEE & JAE  ; 
 FEB <=  KEB & jae  |  KEF & JAE  ; 
 KEB <=  ceb & EEB  |  CEB & eeb  ; 
 KEF <=  cef & EEB  |  CEF & eeb  ; 
 FEC <=  KEC & jae  |  KEG & JAE  ; 
 FED <=  KED & jae  |  KEH & JAE  ; 
 KED <=  ced & EED  |  CED & eed  ; 
 KEH <=  ceh & EED  |  CEH & eed  ; 
 FFA <=  KFA & jaf  |  KFE & JAF  ; 
 FFB <=  KFB & jaf  |  KFF & JAF  ; 
 nae <=  mae & jae  |  mbe & JAE  |  JBB  ; 
 nbe <=  mce & jae  |  mde & JAE  |  jbb  ; 
 UEA <=  SEA & jae  |  SEC & JAE  ; 
 UEB <=  SEB & jae  |  SED & JAE  ; 
 GMC <=  CIE & EJE & EKE & ELE  |  CJE & EKE & ELE  |  CKE & ELE  |  CLE  ; 
 OIA <=  qdb & PAA & PAC & PAB  ; 
 GEA <=  CAE & EBE & ECE & EDE  |  CBE & ECE & EDE  |  CCE & EDE  |  CDE  ; 
 naf <=  maf & jaf  |  mbf & JAF  |  JBA  ; 
 nbf <=  mcf & jaf  |  mdf & JAF  |  jba  ; 
 UFA <=  SFA & jaf  |  SFC & JAF  ; 
 UFB <=  SFB & jaf  |  SFD & JAF  ; 
 KFB <=  cfb & EFB  |  CFB & efb  ; 
 KFF <=  cff & EFB  |  CFF & efb  ; 
 FFC <=  KFC & jaf  |  KFG & JAF  ; 
 FFD <=  KFD & jaf  |  KFH & JAF  ; 
 KFD <=  cfd & EFD  |  CFD & efd  ; 
 KFH <=  cfh & EFD  |  CFH & efd  ; 
 KEA <=  EEA  ; 
 KEE <=  eea  ; 
 ABA <=  IEA & IEA  |  IBA  ; 
 BBA <=  IBA & IEA  ; 
 KEC <=  cec & EEC  |  CEC & eec  ; 
 KEG <=  ceg & EEC  |  CEG & eec  ; 
 ABB <=  IEB & IEB  |  IBB  ; 
 BBB <=  IBB & IEB  ; 
 ABC <=  IEC & IEC  |  IBC  ; 
 BBC <=  IBC & IEC  ; 
 gfa <=  cee & cee  ; 
 gga <=  cfe & cee  |  cfe & efe  ; 
 ABD <=  IED & IED  |  IBD  ; 
 BBD <=  IBD & IED  ; 
 gla <=  ZZO & cie & cje & cke  |  ZZI & cie & cje & cke  |  eje & cje & cke  |  eke & cke & cke  ; 
 ABE <=  IEE & IEE  |  IBE  ; 
 BBE <=  IBE & IEE  ; 
 ABF <=  IEF & IEF  |  IBF  ; 
 BBF <=  IBF & IEF  ; 
 KFA <=  EFA  ; 
 KFE <=  efa  ; 
 ABG <=  IEG & IEG  |  IBG  ; 
 BBG <=  IBG & IEG  ; 
 KFC <=  cfc & EFC  |  CFC & efc  ; 
 KFG <=  cfg & EFC  |  CFG & efc  ; 
 ABH <=  IEH & IEH  |  IBH  ; 
 BBH <=  IBH & IEH  ; 
 FCA <=  KCA & jac  |  KCE & JAC  ; 
 FCB <=  KCB & jac  |  KCF & JAC  ; 
 KCB <=  ccb & ECB  |  CCB & ecb  ; 
 KCF <=  ccf & ECB  |  CCF & ecb  ; 
 FCC <=  KCC & jac  |  KCG & JAC  ; 
 FCD <=  KCD & jac  |  KCH & JAC  ; 
 KCD <=  ccd & ECD  |  CCD & ecd  ; 
 KCH <=  cch & ECD  |  CCH & ecd  ; 
 FDA <=  KDA & jad  |  KDE & JAD  ; 
 FDB <=  KDB & jad  |  KDF & JAD  ; 
 nac <=  mac & jac  |  mbc & JAC  |  JBB  ; 
 nbc <=  mcc & jac  |  mdc & JAC  |  jbb  ; 
 UCA <=  SCA & jac  |  SCC & JAC  ; 
 UCB <=  SCB & jac  |  SCD & JAC  ; 
 GMA <=  CIE & EJE & EKE & ELE  |  CJE & EKE & ELE  |  CKE & ELE  |  CLE  ; 
 nad <=  mad & jad  |  mbd & JAD  |  JBA  ; 
 nbd <=  mcd & jad  |  mdd & JAD  |  jba  ; 
 UDA <=  SDA & jad  |  SDC & JAD  ; 
 UDB <=  SDB & jad  |  SDD & JAD  ; 
 KDB <=  cdb & EDB  |  CDB & edb  ; 
 KDF <=  cdf & EDB  |  CDF & edb  ; 
 FDC <=  KDC & jad  |  KDG & JAD  ; 
 FDD <=  KDD & jad  |  KDH & JAD  ; 
 KDD <=  cdd & EDD  |  CDD & edd  ; 
 KDH <=  cdh & EDD  |  CDH & edd  ; 
 KCA <=  ECA  ; 
 KCE <=  eca  ; 
 gda <=  ZZO & cae & cbe & cce  |  ZZI & cae & cbe & cce  |  ebe & cbe & cce  |  ece & cce & cce  ; 
 AAI <=  IDI & IDI  |  IAI  ; 
 BAI <=  IAI & IDI  ; 
 KCC <=  ccc & ECC  |  CCC & ecc  ; 
 KCG <=  ccg & ECC  |  CCG & ecc  ; 
 AAJ <=  IDJ & IDJ  |  IAJ  ; 
 BAJ <=  IAJ & IDJ  ; 
 AAK <=  IDK & IDK  |  IAK  ; 
 BAK <=  IAK & IDK  ; 
 AAL <=  IDL & IDL  |  IAL  ; 
 BAL <=  IAL & IDL  ; 
 BAO <=  IAO & IDO  ; 
 AAM <=  IDM & IDM  |  IAM  ; 
 BAM <=  IAM & IDM  ; 
 AAN <=  IDN & IDN  |  IAN  ; 
 BAN <=  IAN & IDN  ; 
 KDA <=  EDA  ; 
 KDE <=  eda  ; 
 AAO <=  IDO  |  IAO  ; 
 KDC <=  cdc & EDC  |  CDC & edc  ; 
 KDG <=  cdg & EDC  |  CDG & edc  ; 
 AAP <=  IDP & IDP  |  IAP  ; 
 BAP <=  IAP & IDP  ; 
 FAA <=  KAA & jaa  |  KAE & JAA  ; 
 FAB <=  KAB & jaa  |  KAF & JAA  ; 
 KAB <=  cab & EAB  |  CAB & eab  ; 
 KAF <=  caf & EAB  |  CAF & eab  ; 
 FAC <=  KAC & jaa  |  KAG & JAA  ; 
 FAD <=  KAD & jaa  |  KAH & JAA  ; 
 KAD <=  cad & EAD  |  CAD & ead  ; 
 KAH <=  cah & EAD  |  CAH & ead  ; 
 FBA <=  KBA & jab  |  KBE & JAB  ; 
 FBB <=  KBB & jab  |  KBF & JAB  ; 
 naa <=  maa & jaa  |  mba & JAA  |  JBB  ; 
 UAA <=  SAA & jaa  |  SAC & JAA  ; 
 UAB <=  SAB & jaa  |  SAD & JAA  ; 
 GMB <=  CIE & EJE & EKE & ELE  |  CJE & EKE & ELE  |  CKE & ELE  |  CLE  ; 
 KBB <=  cbb & EBB  |  CBB & ebb  ; 
 ODA <= PAC & PAB ; 
 ODB <= PAC & pab ; 
 nba <=  mca & jaa  |  mda & JAA  |  jbb  ; 
 nab <=  mab & jab  |  mbb & JAB  |  JBA  ; 
 nbb <=  mcb & jab  |  mdb & JAB  |  jba  ; 
 UBA <=  SBA & jab  |  SBC & JAB  ; 
 UBB <=  SBB & jab  |  SBD & JAB  ; 
 KBF <=  cbf & EBB  |  CBF & ebb  ; 
 FBC <=  KBC & jab  |  KBG & JAB  ; 
 FBD <=  KBD & jab  |  KBH & JAB  ; 
 KBD <=  cbd & EBD  |  CBD & ebd  ; 
 KBH <=  cbh & EBD  |  CBH & ebd  ; 
 KAA <= EAA ; 
 KAE <= eaa ; 
 KBA <= EBA ; 
 AAA <=  IAA  |  IDA  |  IAR  ; 
 aar <=  iaa  |  ida  |  iar  ; 
 AAQ <=  IAA & ida & iar  |  iaa & IDA & iar  |  iaa & ida & IAR  |  IAA & IDA & IAR  ;
 baa <=  IAA & ida & iar  |  iaa & IDA & iar  |  iaa & ida & IAR  |  iaa & ida & iar  ;
 KAC <=  cac & EAC  |  CAC & eac  ; 
 KAG <=  cag & EAC  |  CAG & eac  ; 
 FID <=  KID & jai  |  KIH & JAI  ; 
 AAB <=  IDB & IDB  |  IAB  ; 
 BAB <=  IAB & IDB  ; 
 AAC <=  IDC & IDC  |  IAC  ; 
 BAC <=  IAC & IDC  ; 
 gba <=  cae  ; 
 AAD <=  IDD & IDD  |  IAD  ; 
 BAD <=  IAD & IDD  ; 
 hca <=  eie  ; 
 hcb <=  eie  |  eje  ; 
 AAE <=  IDE & IDE  |  IAE  ; 
 BAE <=  IAE & IDE  ; 
 AAF <=  IDF & IDF  |  IAF  ; 
 BAF <=  IAF & IDF  ; 
 KBE <=  eba  ; 
 AAG <=  IDG & IDG  |  IAG  ; 
 BAG <=  IAG & IDG  ; 
 KBC <=  cbc & EBC  |  CBC & ebc  ; 
 KBG <=  cbg & EBC  |  CBG & ebc  ; 
 AAH <=  IDH & IDH  |  IAH  ; 
 BAH <=  IAH & IDH  ; 
 end 
end module
