module bo( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 ICQ, 
 ICR, 
 ICS, 
 ICT, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IGA, 
 IHA, 
 IHB, 
 IHC, 
 IIA, 
 IIB, 
 IIC, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IKI, 
 IKJ, 
 IKK, 
 IKL, 
 ILA, 
 ILB, 
 ILC, 
 ILD, 
 ILE, 
 ILF, 
 ILG, 
 ILH, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 IMH, 
 IXA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OII, 
 OIJ, 
 OIK, 
 OIL, 
 OIM, 
 OIN, 
 OIO, 
 OIP, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OKN, 
 OKO, 
 OKP, 
 OKQ, 
 OKR, 
 OKS, 
 OKT, 
 OLA, 
 OLB, 
 OLC, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 ONA, 
 ONB, 
OOA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input ICQ; 
 input ICR; 
 input ICS; 
 input ICT; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IGA; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IIA; 
 input IIB; 
 input IIC; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IKI; 
 input IKJ; 
 input IKK; 
 input IKL; 
 input ILA; 
 input ILB; 
 input ILC; 
 input ILD; 
 input ILE; 
 input ILF; 
 input ILG; 
 input ILH; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input IMH; 
 input IXA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OII; 
 output OIJ; 
 output OIK; 
 output OIL; 
 output OIM; 
 output OIN; 
 output OIO; 
 output OIP; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OKN; 
 output OKO; 
 output OKP; 
 output OKQ; 
 output OKR; 
 output OKS; 
 output OKT; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output ONA; 
 output ONB; 
 output OOA; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aae ;
reg  aaf ;
reg  aag ;
reg  aah ;
reg  aai ;
reg  aaj ;
reg  aak ;
reg  aal ;
reg  aam ;
reg  aan ;
reg  aao ;
reg  aap ;
reg  aaq ;
reg  aar ;
reg  aas ;
reg  AAT ;
reg  AAU ;
reg  AAV ;
reg  AAW ;
reg  AAX ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  abe ;
reg  abf ;
reg  abg ;
reg  abh ;
reg  abi ;
reg  abj ;
reg  abk ;
reg  abl ;
reg  abm ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  abq ;
reg  abr ;
reg  abs ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  hab ;
reg  hac ;
reg  had ;
reg  hae ;
reg  haf ;
reg  hag ;
reg  hah ;
reg  hai ;
reg  haj ;
reg  hak ;
reg  hal ;
reg  JOA ;
reg  JOB ;
reg  JOC ;
reg  JOD ;
reg  JOE ;
reg  JOF ;
reg  JOG ;
reg  JOH ;
reg  JOI ;
reg  JOJ ;
reg  JOK ;
reg  JOL ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LAG ;
reg  LAH ;
reg  LAI ;
reg  LAJ ;
reg  LAK ;
reg  LAL ;
reg  LAM ;
reg  LAN ;
reg  LAO ;
reg  LAP ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  LBG ;
reg  LBH ;
reg  LBI ;
reg  LBJ ;
reg  LBK ;
reg  LBL ;
reg  LBM ;
reg  LBN ;
reg  LBO ;
reg  LBP ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NCG ;
reg  NCH ;
reg  NCI ;
reg  NCJ ;
reg  NCK ;
reg  NCL ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NDE ;
reg  NDF ;
reg  NDG ;
reg  NDH ;
reg  NDI ;
reg  NDJ ;
reg  NDK ;
reg  NDL ;
reg  NEA ;
reg  NEB ;
reg  NEC ;
reg  NED ;
reg  NEE ;
reg  NEF ;
reg  NEG ;
reg  NEH ;
reg  NEI ;
reg  NEJ ;
reg  NEK ;
reg  NEL ;
reg  NFA ;
reg  NFB ;
reg  NFC ;
reg  NFD ;
reg  NFE ;
reg  NFF ;
reg  NFG ;
reg  NFH ;
reg  NFI ;
reg  NFJ ;
reg  NFK ;
reg  NFL ;
reg  NGA ;
reg  NGB ;
reg  NGC ;
reg  NGD ;
reg  NGE ;
reg  NGF ;
reg  NGG ;
reg  NGH ;
reg  NGI ;
reg  NGJ ;
reg  NGK ;
reg  NGL ;
reg  NHA ;
reg  NHB ;
reg  NHC ;
reg  NHD ;
reg  NHE ;
reg  NHF ;
reg  NHG ;
reg  NHH ;
reg  NHI ;
reg  NHJ ;
reg  NHK ;
reg  NHL ;
reg  NHM ;
reg  NHN ;
reg  NIA ;
reg  NIB ;
reg  NIC ;
reg  NID ;
reg  NIE ;
reg  NIF ;
reg  NIG ;
reg  NIH ;
reg  NII ;
reg  NIJ ;
reg  NIK ;
reg  NIL ;
reg  NIM ;
reg  NIN ;
reg  NJA ;
reg  NJB ;
reg  NJC ;
reg  NJD ;
reg  NJE ;
reg  NJF ;
reg  NJG ;
reg  NJH ;
reg  NJI ;
reg  NJJ ;
reg  NJK ;
reg  NJL ;
reg  NJM ;
reg  NJN ;
reg  NKA ;
reg  NKB ;
reg  NKC ;
reg  NKD ;
reg  NKE ;
reg  NKF ;
reg  NKG ;
reg  NKH ;
reg  NKI ;
reg  NKJ ;
reg  NKK ;
reg  NKL ;
reg  NKM ;
reg  NKN ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  OHL ;
reg  OHM ;
reg  OHN ;
reg  OHO ;
reg  OHP ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OII ;
reg  OIJ ;
reg  OIK ;
reg  OIL ;
reg  OIM ;
reg  OIN ;
reg  OIO ;
reg  OIP ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  ojk ;
reg  ojl ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  OKG ;
reg  OKH ;
reg  OKI ;
reg  OKJ ;
reg  OKK ;
reg  OKL ;
reg  OKM ;
reg  OKN ;
reg  OKO ;
reg  OKP ;
reg  OKQ ;
reg  OKR ;
reg  OKS ;
reg  OKT ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  OME ;
reg  OMF ;
reg  ONA ;
reg  ONB ;
reg  OOA ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  pba ;
reg  pbb ;
reg  pbc ;
reg  pbd ;
reg  pca ;
reg  pcb ;
reg  pcc ;
reg  pcd ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  QAL ;
reg  QAM ;
reg  QAN ;
reg  QAO ;
reg  QAP ;
reg  QAQ ;
reg  QAR ;
reg  QAS ;
reg  QAT ;
reg  QAU ;
reg  QAV ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QBF ;
reg  QBG ;
reg  QBH ;
reg  QBI ;
reg  QBJ ;
reg  QBK ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QEA ;
reg  QEB ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QGA ;
reg  QGB ;
reg  QHA ;
reg  QHB ;
reg  QHC ;
reg  QHD ;
reg  QHE ;
reg  QHF ;
reg  QHG ;
reg  QHH ;
reg  qia ;
reg  QIB ;
reg  qic ;
reg  QID ;
reg  qie ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  qjf ;
reg  QJG ;
reg  QJH ;
reg  QJI ;
reg  QJJ ;
reg  qjo ;
reg  qjp ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  qlf ;
reg  qlg ;
reg  QLH ;
reg  QLI ;
reg  QLJ ;
reg  QLK ;
reg  qll ;
reg  QMA ;
reg  QMB ;
reg  QMC ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  qoa ;
reg  QOB ;
reg  QOC ;
reg  QOD ;
reg  QOF ;
reg  QPA ;
reg  QPB ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  qsa ;
reg  qsb ;
reg  qsc ;
reg  qsd ;
reg  QSE ;
reg  QTB ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QUD ;
reg  QUE ;
reg  QUF ;
reg  QUG ;
reg  QUH ;
reg  QUI ;
reg  QUJ ;
reg  QUK ;
reg  QUL ;
reg  QUM ;
reg  QUN ;
reg  QVD ;
reg  QVE ;
reg  QVF ;
reg  QVG ;
reg  QVH ;
reg  QVI ;
reg  QVJ ;
reg  QVK ;
reg  QWA ;
reg  QWB ;
reg  QWC ;
reg  QWD ;
reg  QWE ;
reg  QWF ;
reg  QWG ;
reg  QWH ;
reg  QXA ;
reg  QXB ;
reg  QXC ;
reg  QXD ;
reg  QXE ;
reg  QXF ;
reg  QXG ;
reg  QXH ;
reg  QZA ;
reg  QZB ;
reg  QZC ;
reg  QZD ;
reg  QZE ;
reg  QZF ;
reg  QZG ;
reg  QZH ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  SAD ;
reg  SAE ;
reg  SAF ;
reg  SAG ;
reg  SAH ;
reg  SAI ;
reg  SAJ ;
reg  SAK ;
reg  SAL ;
reg  SAM ;
reg  SAN ;
reg  SAO ;
reg  SAP ;
reg  SAQ ;
reg  SAR ;
reg  SAS ;
reg  SAT ;
reg  SAU ;
reg  SAV ;
reg  SAW ;
reg  SAX ;
reg  SBA ;
reg  SBB ;
reg  SBC ;
reg  SCA ;
reg  SCB ;
reg  SCC ;
reg  SCD ;
reg  SCE ;
reg  SCF ;
reg  SCG ;
reg  SCH ;
reg  SCI ;
reg  SCJ ;
reg  SCK ;
reg  SCL ;
reg  SDM ;
reg  SEM ;
reg  SFM ;
reg  tbb ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
reg  tga ;
reg  tgb ;
reg  tgc ;
reg  tgd ;
reg  THA ;
reg  THB ;
reg  THC ;
reg  THD ;
reg  THE ;
reg  THF ;
reg  THG ;
reg  THH ;
reg  THI ;
reg  THJ ;
reg  THK ;
reg  THL ;
reg  TIA ;
reg  TIB ;
reg  VAA ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WEA ;
reg  WEB ;
reg  WEC ;
reg  WED ;
reg  WFA ;
reg  WFB ;
reg  WFC ;
reg  WFD ;
reg  WGA ;
reg  WGB ;
reg  WGC ;
reg  WGD ;
reg  WHA ;
reg  WHB ;
reg  WHC ;
reg  WHD ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  AAE ;
wire  AAF ;
wire  AAG ;
wire  AAH ;
wire  AAI ;
wire  AAJ ;
wire  AAK ;
wire  AAL ;
wire  AAM ;
wire  AAN ;
wire  AAO ;
wire  AAP ;
wire  AAQ ;
wire  AAR ;
wire  AAS ;
wire  aat ;
wire  aau ;
wire  aav ;
wire  aaw ;
wire  aax ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ABE ;
wire  ABF ;
wire  ABG ;
wire  ABH ;
wire  ABI ;
wire  ABJ ;
wire  ABK ;
wire  ABL ;
wire  ABM ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  ABQ ;
wire  ABR ;
wire  ABS ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fam ;
wire  FAM ;
wire  fan ;
wire  FAN ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  fbi ;
wire  FBI ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbl ;
wire  FBL ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fcg ;
wire  FCG ;
wire  fch ;
wire  FCH ;
wire  fci ;
wire  FCI ;
wire  fcj ;
wire  FCJ ;
wire  fck ;
wire  FCK ;
wire  fcl ;
wire  FCL ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fdh ;
wire  FDH ;
wire  fdi ;
wire  FDI ;
wire  fdj ;
wire  FDJ ;
wire  fdk ;
wire  FDK ;
wire  fdl ;
wire  FDL ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gai ;
wire  GAI ;
wire  gaj ;
wire  GAJ ;
wire  gak ;
wire  GAK ;
wire  gal ;
wire  GAL ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  HAE ;
wire  HAF ;
wire  HAG ;
wire  HAH ;
wire  HAI ;
wire  HAJ ;
wire  HAK ;
wire  HAL ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  icq ;
wire  icr ;
wire  ics ;
wire  ict ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  iga ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  iia ;
wire  iib ;
wire  iic ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  iki ;
wire  ikj ;
wire  ikk ;
wire  ikl ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ild ;
wire  ile ;
wire  ilf ;
wire  ilg ;
wire  ilh ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  imh ;
wire  ixa ;
wire  jaa ;
wire  JAA ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jga ;
wire  JGA ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  jne ;
wire  JNE ;
wire  jnf ;
wire  JNF ;
wire  joa ;
wire  job ;
wire  joc ;
wire  jod ;
wire  joe ;
wire  jof ;
wire  jog ;
wire  joh ;
wire  joi ;
wire  joj ;
wire  jok ;
wire  jol ;
wire  jpa ;
wire  JPA ;
wire  jpb ;
wire  JPB ;
wire  jpc ;
wire  JPC ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lag ;
wire  lah ;
wire  lai ;
wire  laj ;
wire  lak ;
wire  lal ;
wire  lam ;
wire  lan ;
wire  lao ;
wire  lap ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  lbg ;
wire  lbh ;
wire  lbi ;
wire  lbj ;
wire  lbk ;
wire  lbl ;
wire  lbm ;
wire  lbn ;
wire  lbo ;
wire  lbp ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  ncg ;
wire  nch ;
wire  nci ;
wire  ncj ;
wire  nck ;
wire  ncl ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nde ;
wire  ndf ;
wire  ndg ;
wire  ndh ;
wire  ndi ;
wire  ndj ;
wire  ndk ;
wire  ndl ;
wire  nea ;
wire  neb ;
wire  nec ;
wire  ned ;
wire  nee ;
wire  nef ;
wire  neg ;
wire  neh ;
wire  nei ;
wire  nej ;
wire  nek ;
wire  nel ;
wire  nfa ;
wire  nfb ;
wire  nfc ;
wire  nfd ;
wire  nfe ;
wire  nff ;
wire  nfg ;
wire  nfh ;
wire  nfi ;
wire  nfj ;
wire  nfk ;
wire  nfl ;
wire  nga ;
wire  ngb ;
wire  ngc ;
wire  ngd ;
wire  nge ;
wire  ngf ;
wire  ngg ;
wire  ngh ;
wire  ngi ;
wire  ngj ;
wire  ngk ;
wire  ngl ;
wire  nha ;
wire  nhb ;
wire  nhc ;
wire  nhd ;
wire  nhe ;
wire  nhf ;
wire  nhg ;
wire  nhh ;
wire  nhi ;
wire  nhj ;
wire  nhk ;
wire  nhl ;
wire  nhm ;
wire  nhn ;
wire  nia ;
wire  nib ;
wire  nic ;
wire  nid ;
wire  nie ;
wire  nif ;
wire  nig ;
wire  nih ;
wire  nii ;
wire  nij ;
wire  nik ;
wire  nil ;
wire  nim ;
wire  nin ;
wire  nja ;
wire  njb ;
wire  njc ;
wire  njd ;
wire  nje ;
wire  njf ;
wire  njg ;
wire  njh ;
wire  nji ;
wire  njj ;
wire  njk ;
wire  njl ;
wire  njm ;
wire  njn ;
wire  nka ;
wire  nkb ;
wire  nkc ;
wire  nkd ;
wire  nke ;
wire  nkf ;
wire  nkg ;
wire  nkh ;
wire  nki ;
wire  nkj ;
wire  nkk ;
wire  nkl ;
wire  nkm ;
wire  nkn ;
wire  nla ;
wire  NLA ;
wire  nlb ;
wire  NLB ;
wire  nlc ;
wire  NLC ;
wire  nld ;
wire  NLD ;
wire  nle ;
wire  NLE ;
wire  nlf ;
wire  NLF ;
wire  nlg ;
wire  NLG ;
wire  nlh ;
wire  NLH ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  ohl ;
wire  ohm ;
wire  ohn ;
wire  oho ;
wire  ohp ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oii ;
wire  oij ;
wire  oik ;
wire  oil ;
wire  oim ;
wire  oin ;
wire  oio ;
wire  oip ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  OJK ;
wire  OJL ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  okg ;
wire  okh ;
wire  oki ;
wire  okj ;
wire  okk ;
wire  okl ;
wire  okm ;
wire  okn ;
wire  oko ;
wire  okp ;
wire  okq ;
wire  okr ;
wire  oks ;
wire  okt ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  ome ;
wire  omf ;
wire  ona ;
wire  onb ;
wire  ooa ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  PBA ;
wire  PBB ;
wire  PBC ;
wire  PBD ;
wire  PCA ;
wire  PCB ;
wire  PCC ;
wire  PCD ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  qal ;
wire  qam ;
wire  qan ;
wire  qao ;
wire  qap ;
wire  qaq ;
wire  qar ;
wire  qas ;
wire  qat ;
wire  qau ;
wire  qav ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qbf ;
wire  qbg ;
wire  qbh ;
wire  qbi ;
wire  qbj ;
wire  qbk ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qea ;
wire  qeb ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qga ;
wire  qgb ;
wire  qha ;
wire  qhb ;
wire  qhc ;
wire  qhd ;
wire  qhe ;
wire  qhf ;
wire  qhg ;
wire  qhh ;
wire  QIA ;
wire  qib ;
wire  QIC ;
wire  qid ;
wire  QIE ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  QJF ;
wire  qjg ;
wire  qjh ;
wire  qji ;
wire  qjj ;
wire  qjk ;
wire  QJK ;
wire  qjl ;
wire  QJL ;
wire  qjm ;
wire  QJM ;
wire  qjn ;
wire  QJN ;
wire  QJO ;
wire  QJP ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  QLF ;
wire  QLG ;
wire  qlh ;
wire  qli ;
wire  qlj ;
wire  qlk ;
wire  QLL ;
wire  qma ;
wire  qmb ;
wire  qmc ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  QOA ;
wire  qob ;
wire  qoc ;
wire  qod ;
wire  qof ;
wire  qpa ;
wire  qpb ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  QSA ;
wire  QSB ;
wire  QSC ;
wire  QSD ;
wire  qse ;
wire  qtb ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qud ;
wire  que ;
wire  quf ;
wire  qug ;
wire  quh ;
wire  qui ;
wire  quj ;
wire  quk ;
wire  qul ;
wire  qum ;
wire  qun ;
wire  qvd ;
wire  qve ;
wire  qvf ;
wire  qvg ;
wire  qvh ;
wire  qvi ;
wire  qvj ;
wire  qvk ;
wire  qwa ;
wire  qwb ;
wire  qwc ;
wire  qwd ;
wire  qwe ;
wire  qwf ;
wire  qwg ;
wire  qwh ;
wire  qxa ;
wire  qxb ;
wire  qxc ;
wire  qxd ;
wire  qxe ;
wire  qxf ;
wire  qxg ;
wire  qxh ;
wire  qya ;
wire  QYA ;
wire  qyb ;
wire  QYB ;
wire  qza ;
wire  qzb ;
wire  qzc ;
wire  qzd ;
wire  qze ;
wire  qzf ;
wire  qzg ;
wire  qzh ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  saa ;
wire  sab ;
wire  sac ;
wire  sad ;
wire  sae ;
wire  saf ;
wire  sag ;
wire  sah ;
wire  sai ;
wire  saj ;
wire  sak ;
wire  sal ;
wire  sam ;
wire  san ;
wire  sao ;
wire  sap ;
wire  saq ;
wire  sar ;
wire  sas ;
wire  sat ;
wire  sau ;
wire  sav ;
wire  saw ;
wire  sax ;
wire  sba ;
wire  sbb ;
wire  sbc ;
wire  sca ;
wire  scb ;
wire  scc ;
wire  scd ;
wire  sce ;
wire  scf ;
wire  scg ;
wire  sch ;
wire  sci ;
wire  scj ;
wire  sck ;
wire  scl ;
wire  sdm ;
wire  sem ;
wire  sfm ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tae ;
wire  TAE ;
wire  taf ;
wire  TAF ;
wire  tag ;
wire  TAG ;
wire  tah ;
wire  TAH ;
wire  tai ;
wire  TAI ;
wire  taj ;
wire  TAJ ;
wire  tba ;
wire  TBA ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tbe ;
wire  TBE ;
wire  tbf ;
wire  TBF ;
wire  tbg ;
wire  TBG ;
wire  tbh ;
wire  TBH ;
wire  tbi ;
wire  TBI ;
wire  tbm ;
wire  TBM ;
wire  tbn ;
wire  TBN ;
wire  tbo ;
wire  TBO ;
wire  tbp ;
wire  TBP ;
wire  tbq ;
wire  TBQ ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tda ;
wire  TDA ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  TGA ;
wire  TGB ;
wire  TGC ;
wire  TGD ;
wire  tha ;
wire  thb ;
wire  thc ;
wire  thd ;
wire  the ;
wire  thf ;
wire  thg ;
wire  thh ;
wire  thi ;
wire  thj ;
wire  thk ;
wire  thl ;
wire  tia ;
wire  tib ;
wire  vaa ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wea ;
wire  web ;
wire  wec ;
wire  wed ;
wire  wfa ;
wire  wfb ;
wire  wfc ;
wire  wfd ;
wire  wga ;
wire  wgb ;
wire  wgc ;
wire  wgd ;
wire  wha ;
wire  whb ;
wire  whc ;
wire  whd ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign saa = ~SAA;  //complement 
assign nka = ~NKA;  //complement 
assign sai = ~SAI;  //complement 
assign nki = ~NKI;  //complement 
assign qau = ~QAU;  //complement 
assign qav = ~QAV;  //complement 
assign saq = ~SAQ;  //complement 
assign raa = ~RAA;  //complement 
assign qla = ~QLA;  //complement 
assign tca =  qaj & qhc  ; 
assign TCA = ~tca;  //complement 
assign qlb = ~QLB;  //complement 
assign qad = ~QAD;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign qai = ~QAI;  //complement 
assign qaj = ~QAJ;  //complement 
assign qak = ~QAK;  //complement 
assign qal = ~QAL;  //complement 
assign qam = ~QAM;  //complement 
assign qan = ~QAN;  //complement 
assign qao = ~QAO;  //complement 
assign qap = ~QAP;  //complement 
assign qaq = ~QAQ;  //complement 
assign sba = ~SBA;  //complement 
assign omf = ~OMF;  //complement 
assign kaa = ~KAA;  //complement 
assign kai = ~KAI;  //complement 
assign oka = ~OKA;  //complement 
assign baa = ~BAA;  //complement 
assign bai = ~BAI;  //complement 
assign TAA = qia & qob ; 
assign taa = ~TAA ; //complement 
assign TAJ = qia & qob ; 
assign taj = ~TAJ ;  //complement 
assign tad = qia & ZZI ; 
assign TAD = ~tad ;  //complement 
assign oia = ~OIA;  //complement 
assign oii = ~OII;  //complement 
assign AAA = ~aaa;  //complement 
assign AAI = ~aai;  //complement 
assign ABA = ~aba;  //complement 
assign ABI = ~abi;  //complement 
assign QIA = ~qia;  //complement 
assign QIE = ~qie;  //complement 
assign daa = ~DAA;  //complement 
assign OJK = ~ojk;  //complement 
assign OJL = ~ojl;  //complement 
assign aat = ~AAT;  //complement 
assign oha = ~OHA;  //complement 
assign ohi = ~OHI;  //complement 
assign oki = ~OKI;  //complement 
assign qaa = ~QAA;  //complement 
assign JBA =  aal & aak & aaj  ; 
assign jba = ~JBA;  //complement 
assign tda =  qaa & qca  ; 
assign TDA = ~tda;  //complement 
assign NLA =  RAA & QLK  ; 
assign nla = ~NLA;  //complement 
assign jma = abq & qma ; 
assign JMA = ~jma ; //complement 
assign jmb = abq & qma ; 
assign JMB = ~jmb ;  //complement 
assign okq = ~OKQ;  //complement 
assign QIC = ~qic;  //complement 
assign qma = ~QMA;  //complement 
assign olc = ~OLC;  //complement 
assign qab = ~QAB;  //complement 
assign qob = ~QOB;  //complement 
assign qof = ~QOF;  //complement 
assign omb = ~OMB;  //complement 
assign AAQ = ~aaq;  //complement 
assign ABQ = ~abq;  //complement 
assign omc = ~OMC;  //complement 
assign omd = ~OMD;  //complement 
assign qac = ~QAC;  //complement 
assign qas = ~QAS;  //complement 
assign JGA =  QLA & qib  |  QLB & qib  ; 
assign jga = ~JGA;  //complement 
assign qar = ~QAR;  //complement 
assign qib = ~QIB;  //complement 
assign gaa =  NDA & ZZI & QNA  |  ZZI & ZZO  |  naa & qna  ; 
assign GAA = ~gaa; //complement 
assign gad =  NDD & HAD & QNA  |  nad & had  |  nad & qna  ; 
assign GAD = ~gad; //complement 
assign gag =  NDG & HAG & QNB  |  nag & hag  |  nag & qnb  ; 
assign GAG = ~gag; //complement 
assign gaj =  NDJ & HAJ & QNC  |  naj & haj  |  naj & qnc  ; 
assign GAJ = ~gaj; //complement 
assign HAD = ~had;  //complement 
assign HAG = ~hag;  //complement 
assign HAJ = ~haj;  //complement 
assign sab = ~SAB;  //complement 
assign nkb = ~NKB;  //complement 
assign saj = ~SAJ;  //complement 
assign nkj = ~NKJ;  //complement 
assign sar = ~SAR;  //complement 
assign rab = ~RAB;  //complement 
assign tcb =  qaj & qhc  ; 
assign TCB = ~tcb;  //complement 
assign jda =  qbd & qbg & qbh  ; 
assign JDA = ~jda;  //complement 
assign qlc = ~QLC;  //complement 
assign qld = ~QLD;  //complement 
assign qbb = ~QBB;  //complement 
assign qbc = ~QBC;  //complement 
assign qbd = ~QBD;  //complement 
assign qbe = ~QBE;  //complement 
assign qbf = ~QBF;  //complement 
assign qbg = ~QBG;  //complement 
assign qbh = ~QBH;  //complement 
assign qbi = ~QBI;  //complement 
assign tbf =  qlc  ; 
assign TBF = ~tbf;  //complement 
assign tba =  qlc  ; 
assign TBA = ~tba;  //complement 
assign tbp =  qlc  ; 
assign TBP = ~tbp;  //complement 
assign kab = ~KAB;  //complement 
assign kaj = ~KAJ;  //complement 
assign okb = ~OKB;  //complement 
assign bab = ~BAB;  //complement 
assign baj = ~BAJ;  //complement 
assign TAB = QLC; 
assign tab = ~TAB; //complement 
assign tah = qia; 
assign TAH = ~tah;  //complement 
assign TAE = qie & qof ; 
assign tae = ~TAE ;  //complement 
assign TAI = qie & qob; 
assign tai = ~TAI; 
assign oib = ~OIB;  //complement 
assign oij = ~OIJ;  //complement 
assign AAB = ~aab;  //complement 
assign AAJ = ~aaj;  //complement 
assign ABB = ~abb;  //complement 
assign aau = ~AAU;  //complement 
assign TAF = QLC; 
assign taf = ~TAF; //complement 
assign TAC = QLD; 
assign tac = ~TAC;  //complement 
assign TAG = QLD; 
assign tag = ~TAG;  //complement 
assign dab = ~DAB;  //complement 
assign qje = ~QJE;  //complement 
assign QOA = ~qoa;  //complement 
assign acj = ~ACJ;  //complement 
assign ohb = ~OHB;  //complement 
assign ohj = ~OHJ;  //complement 
assign okj = ~OKJ;  //complement 
assign qba = ~QBA;  //complement 
assign JBB =  aal & aak & AAU  ; 
assign jbb = ~JBB;  //complement 
assign NLB =  RAB & QLK  ; 
assign nlb = ~NLB;  //complement 
assign JAA =  ABR & aap & aao & aan & AAX  ; 
assign jaa = ~JAA;  //complement  
assign okr = ~OKR;  //complement 
assign sbb = ~SBB;  //complement 
assign qbj = ~QBJ;  //complement 
assign qjc = ~QJC;  //complement 
assign AAR = ~aar;  //complement 
assign ABR = ~abr;  //complement 
assign ABJ = ~abj;  //complement 
assign qbk = ~QBK;  //complement 
assign qtb = ~QTB;  //complement 
assign quc = ~QUC;  //complement 
assign qud = ~QUD;  //complement 
assign que = ~QUE;  //complement 
assign quf = ~QUF;  //complement 
assign qua = ~QUA;  //complement 
assign qub = ~QUB;  //complement 
assign QSA = ~qsa;  //complement 
assign QSB = ~qsb;  //complement 
assign QSC = ~qsc;  //complement 
assign QSD = ~qsd;  //complement 
assign gab =  NDB & HAB & QNA  |  nab & hab  |  nab & qna  ; 
assign GAB = ~gab; //complement 
assign gae =  NDE & HAE & QNB  |  nae & hae  |  nae & qnb  ; 
assign GAE = ~gae; //complement 
assign gah =  NDH & HAH & QNB  |  nah & hah  |  nah & qnb  ; 
assign GAH = ~gah; //complement 
assign gak =  NDK & HAK & QNC  |  nak & hak  |  nak & qnc  ; 
assign GAK = ~gak; //complement 
assign HAB = ~hab;  //complement 
assign HAE = ~hae;  //complement 
assign HAH = ~hah;  //complement 
assign HAK = ~hak;  //complement 
assign sac = ~SAC;  //complement 
assign nkc = ~NKC;  //complement 
assign qpa = ~QPA;  //complement 
assign qpb = ~QPB;  //complement 
assign sak = ~SAK;  //complement 
assign nkk = ~NKK;  //complement 
assign qra = ~QRA;  //complement 
assign qrb = ~QRB;  //complement 
assign qrc = ~QRC;  //complement 
assign qse = ~QSE;  //complement 
assign sas = ~SAS;  //complement 
assign rac = ~RAC;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tec = ~TEC;  //complement 
assign ted = ~TED;  //complement 
assign qrd = ~QRD;  //complement 
assign qre = ~QRE;  //complement 
assign tcc =  qaj & qhc  ; 
assign TCC = ~tcc;  //complement 
assign tcd =  qat & qhd  ; 
assign TCD = ~tcd;  //complement 
assign tce =  qat & qhd  ; 
assign TCE = ~tce;  //complement 
assign qhc = ~QHC;  //complement 
assign qhd = ~QHD;  //complement 
assign qat = ~QAT;  //complement 
assign qhe = ~QHE;  //complement 
assign qhf = ~QHF;  //complement 
assign qhg = ~QHG;  //complement 
assign qhh = ~QHH;  //complement 
assign tbq =  qlg  ; 
assign TBQ = ~tbq;  //complement 
assign kac = ~KAC;  //complement 
assign kak = ~KAK;  //complement 
assign okc = ~OKC;  //complement 
assign bac = ~BAC;  //complement 
assign bak = ~BAK;  //complement 
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign oic = ~OIC;  //complement 
assign oik = ~OIK;  //complement 
assign AAC = ~aac;  //complement 
assign AAK = ~aak;  //complement 
assign ABC = ~abc;  //complement 
assign aav = ~AAV;  //complement 
assign sbc = ~SBC;  //complement 
assign dac = ~DAC;  //complement 
assign qjd = ~QJD;  //complement 
assign ack = ~ACK;  //complement 
assign ABK = ~abk;  //complement 
assign ohc = ~OHC;  //complement 
assign ohk = ~OHK;  //complement 
assign okk = ~OKK;  //complement 
assign qca = ~QCA;  //complement 
assign JBC =  aal & AAV & aaj  ; 
assign jbc = ~JBC;  //complement 
assign NLC =  RAC & QLK  ; 
assign nlc = ~NLC;  //complement 
assign qjg = ~QJG;  //complement 
assign qjh = ~QJH;  //complement 
assign qji = ~QJI;  //complement 
assign qjj = ~QJJ;  //complement 
assign oks = ~OKS;  //complement 
assign qcb = ~QCB;  //complement 
assign AAS = ~aas;  //complement 
assign qqa = ~QQA;  //complement 
assign qqb = ~QQB;  //complement 
assign qqc = ~QQC;  //complement 
assign qcc = ~QCC;  //complement 
assign ABS = ~abs;  //complement 
assign ome = ~OME;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign gac =  NDC & HAC & QNA  |  nac & hac  |  nac & qna  ; 
assign GAC = ~gac; //complement 
assign gaf =  NDF & HAF & QNB  |  naf & haf  |  naf & qnb  ; 
assign GAF = ~gaf; //complement 
assign gai =  NDI & HAI & QNC  |  nai & hai  |  nai & qnc  ; 
assign GAI = ~gai; //complement 
assign gal =  NDL & HAL & QNC  |  nal & hal  |  nal & qnc  ; 
assign GAL = ~gal; //complement 
assign HAC = ~hac;  //complement 
assign HAF = ~haf;  //complement 
assign HAI = ~hai;  //complement 
assign HAL = ~hal;  //complement 
assign paa = ~PAA;  //complement 
assign pab = ~PAB;  //complement 
assign pac = ~PAC;  //complement 
assign pad = ~PAD;  //complement 
assign PBA = ~pba;  //complement 
assign PCA = ~pca;  //complement 
assign PBB = ~pbb;  //complement 
assign PCB = ~pcb;  //complement 
assign PBC = ~pbc;  //complement 
assign PCC = ~pcc;  //complement 
assign PBD = ~pbd;  //complement 
assign PCD = ~pcd;  //complement 
assign sad = ~SAD;  //complement 
assign nkd = ~NKD;  //complement 
assign sal = ~SAL;  //complement 
assign nkl = ~NKL;  //complement 
assign sat = ~SAT;  //complement 
assign rad = ~RAD;  //complement 
assign qna = ~QNA;  //complement 
assign qnb = ~QNB;  //complement 
assign qnc = ~QNC;  //complement 
assign lbm = ~LBM;  //complement 
assign lbn = ~LBN;  //complement 
assign lbo = ~LBO;  //complement 
assign lbp = ~LBP;  //complement 
assign qdd = ~QDD;  //complement 
assign tbd =  qll  ; 
assign TBD = ~tbd;  //complement 
assign TBB = ~tbb;  //complement 
assign kal = ~KAL;  //complement 
assign kam = ~KAM;  //complement 
assign okd = ~OKD;  //complement 
assign bad = ~BAD;  //complement 
assign bal = ~BAL;  //complement 
assign kad = ~KAD;  //complement 
assign oid = ~OID;  //complement 
assign oil = ~OIL;  //complement 
assign AAD = ~aad;  //complement 
assign AAL = ~aal;  //complement 
assign ABD = ~abd;  //complement 
assign aaw = ~AAW;  //complement 
assign dad = ~DAD;  //complement 
assign qod = ~QOD;  //complement 
assign acl = ~ACL;  //complement 
assign ABL = ~abl;  //complement 
assign ohd = ~OHD;  //complement 
assign ohl = ~OHL;  //complement 
assign okl = ~OKL;  //complement 
assign qda = ~QDA;  //complement 
assign JBD =  aal & AAV & AAU  ; 
assign jbd = ~JBD;  //complement 
assign NLD =  RAD & QLK  ; 
assign nld = ~NLD;  //complement 
assign jcf =  qaa & qbk & qcc & qdc & qea & qfb  ; 
assign JCF = ~jcf;  //complement  
assign jcg =  qga & qha  ; 
assign JCG = ~jcg;  //complement 
assign okt = ~OKT;  //complement 
assign qoc = ~QOC;  //complement 
assign qdb = ~QDB;  //complement 
assign oma = ~OMA;  //complement 
assign qdc = ~QDC;  //complement 
assign lam = ~LAM;  //complement 
assign lan = ~LAN;  //complement 
assign lao = ~LAO;  //complement 
assign lap = ~LAP;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign thc = ~THC;  //complement 
assign thd = ~THD;  //complement 
assign qvd = ~QVD;  //complement 
assign the = ~THE;  //complement 
assign thf = ~THF;  //complement 
assign thg = ~THG;  //complement 
assign thh = ~THH;  //complement 
assign nad = ~NAD;  //complement 
assign nae = ~NAE;  //complement 
assign naf = ~NAF;  //complement 
assign vaa = ~VAA;  //complement 
assign TGA = ~tga;  //complement 
assign waa = ~WAA;  //complement 
assign wba = ~WBA;  //complement 
assign wca = ~WCA;  //complement 
assign naa = ~NAA;  //complement 
assign nab = ~NAB;  //complement 
assign nac = ~NAC;  //complement 
assign nag = ~NAG;  //complement 
assign nah = ~NAH;  //complement 
assign nai = ~NAI;  //complement 
assign naj = ~NAJ;  //complement 
assign nak = ~NAK;  //complement 
assign nal = ~NAL;  //complement 
assign faa = naa; 
assign FAA = ~faa; //complement 
assign fab = nab; 
assign FAB = ~fab;  //complement 
assign fac = nac; 
assign FAC = ~fac;  //complement 
assign fan = nae; 
assign FAN = ~fan;  //complement 
assign fad = nad; 
assign FAD = ~fad; //complement 
assign fam = nad; 
assign FAM = ~fam;  //complement 
assign fae = nae; 
assign FAE = ~fae;  //complement 
assign faf = naf; 
assign FAF = ~faf;  //complement 
assign wda = ~WDA;  //complement 
assign wea = ~WEA;  //complement 
assign wfa = ~WFA;  //complement 
assign fag =  nag  ; 
assign FAG = ~fag;  //complement 
assign fah =  nah  ; 
assign FAH = ~fah;  //complement 
assign fai =  nai  ; 
assign FAI = ~fai;  //complement 
assign faj =  naj  ; 
assign FAJ = ~faj;  //complement 
assign fak =  nak  ; 
assign FAK = ~fak;  //complement 
assign fal =  nal  ; 
assign FAL = ~fal;  //complement 
assign wga = ~WGA;  //complement 
assign wha = ~WHA;  //complement 
assign JNA =  NAA & NAB & NAC  ; 
assign jna = ~JNA;  //complement 
assign JNB =  NAA & NAB & NAC  ; 
assign jnb = ~JNB;  //complement 
assign JNC =  NAA & NAB & NAC  ; 
assign jnc = ~JNC;  //complement 
assign JND =  NAD & NAE & NAF  ; 
assign jnd = ~JND;  //complement 
assign JNE =  NAD & NAE & NAF  ; 
assign jne = ~JNE;  //complement 
assign JNF =  NAG & NAH & NAI  ; 
assign jnf = ~JNF;  //complement 
assign nea = ~NEA;  //complement 
assign neb = ~NEB;  //complement 
assign nec = ~NEC;  //complement 
assign ned = ~NED;  //complement 
assign nee = ~NEE;  //complement 
assign nef = ~NEF;  //complement 
assign neg = ~NEG;  //complement 
assign neh = ~NEH;  //complement 
assign nei = ~NEI;  //complement 
assign nej = ~NEJ;  //complement 
assign nek = ~NEK;  //complement 
assign nel = ~NEL;  //complement 
assign nfa = ~NFA;  //complement 
assign nfb = ~NFB;  //complement 
assign nfc = ~NFC;  //complement 
assign nfd = ~NFD;  //complement 
assign nhm = ~NHM;  //complement 
assign nhn = ~NHN;  //complement 
assign sae = ~SAE;  //complement 
assign nke = ~NKE;  //complement 
assign JPA =  QRD  ; 
assign jpa = ~JPA;  //complement 
assign jqa =  qau & qmc  ; 
assign JQA = ~jqa;  //complement 
assign JRA =  QAV  ; 
assign jra = ~JRA;  //complement 
assign sam = ~SAM;  //complement 
assign sdm = ~SDM;  //complement 
assign sem = ~SEM;  //complement 
assign nkm = ~NKM;  //complement 
assign lba = ~LBA;  //complement 
assign lbb = ~LBB;  //complement 
assign lbc = ~LBC;  //complement 
assign lbd = ~LBD;  //complement 
assign sau = ~SAU;  //complement 
assign rae = ~RAE;  //complement 
assign sca = ~SCA;  //complement 
assign scb = ~SCB;  //complement 
assign joa = ~JOA;  //complement 
assign job = ~JOB;  //complement 
assign joc = ~JOC;  //complement 
assign jod = ~JOD;  //complement 
assign qeb = ~QEB;  //complement 
assign scc = ~SCC;  //complement 
assign scd = ~SCD;  //complement 
assign nhe = ~NHE;  //complement 
assign nhf = ~NHF;  //complement 
assign nhg = ~NHG;  //complement 
assign nhh = ~NHH;  //complement 
assign nia = ~NIA;  //complement 
assign nib = ~NIB;  //complement 
assign nic = ~NIC;  //complement 
assign nid = ~NID;  //complement 
assign nga = ~NGA;  //complement 
assign ngb = ~NGB;  //complement 
assign ngc = ~NGC;  //complement 
assign ngd = ~NGD;  //complement 
assign nge = ~NGE;  //complement 
assign ngf = ~NGF;  //complement 
assign ngg = ~NGG;  //complement 
assign ngh = ~NGH;  //complement 
assign nie = ~NIE;  //complement 
assign nif = ~NIF;  //complement 
assign nig = ~NIG;  //complement 
assign nih = ~NIH;  //complement 
assign nfi = ~NFI;  //complement 
assign nfj = ~NFJ;  //complement 
assign nfk = ~NFK;  //complement 
assign nfl = ~NFL;  //complement 
assign ngi = ~NGI;  //complement 
assign ngj = ~NGJ;  //complement 
assign ngk = ~NGK;  //complement 
assign ngl = ~NGL;  //complement 
assign nii = ~NII;  //complement 
assign nij = ~NIJ;  //complement 
assign nik = ~NIK;  //complement 
assign nil = ~NIL;  //complement 
assign nfe = ~NFE;  //complement 
assign nff = ~NFF;  //complement 
assign nfg = ~NFG;  //complement 
assign nfh = ~NFH;  //complement 
assign nhi = ~NHI;  //complement 
assign nhj = ~NHJ;  //complement 
assign nhk = ~NHK;  //complement 
assign nhl = ~NHL;  //complement 
assign kae = ~KAE;  //complement 
assign eam =  aam  ; 
assign EAM = ~eam;  //complement 
assign oke = ~OKE;  //complement 
assign bae = ~BAE;  //complement 
assign bam = ~BAM;  //complement 
assign sfm = ~SFM;  //complement 
assign oie = ~OIE;  //complement 
assign oim = ~OIM;  //complement 
assign AAE = ~aae;  //complement 
assign AAM = ~aam;  //complement 
assign ABE = ~abe;  //complement 
assign aax = ~AAX;  //complement 
assign nha = ~NHA;  //complement 
assign nhb = ~NHB;  //complement 
assign nhc = ~NHC;  //complement 
assign nhd = ~NHD;  //complement 
assign dae = ~DAE;  //complement 
assign ABM = ~abm;  //complement 
assign ohe = ~OHE;  //complement 
assign ohm = ~OHM;  //complement 
assign okm = ~OKM;  //complement 
assign qea = ~QEA;  //complement 
assign JBE =  AAW & aak & aaj  ; 
assign jbe = ~JBE;  //complement 
assign NLE =  RAE & QLJ  ; 
assign nle = ~NLE;  //complement 
assign laa = ~LAA;  //complement 
assign lab = ~LAB;  //complement 
assign lac = ~LAC;  //complement 
assign lad = ~LAD;  //complement 
assign nja = ~NJA;  //complement 
assign njb = ~NJB;  //complement 
assign njc = ~NJC;  //complement 
assign njd = ~NJD;  //complement 
assign nje = ~NJE;  //complement 
assign njf = ~NJF;  //complement 
assign njg = ~NJG;  //complement 
assign njh = ~NJH;  //complement 
assign nji = ~NJI;  //complement 
assign njj = ~NJJ;  //complement 
assign njk = ~NJK;  //complement 
assign njl = ~NJL;  //complement 
assign nim = ~NIM;  //complement 
assign nin = ~NIN;  //complement 
assign njm = ~NJM;  //complement 
assign njn = ~NJN;  //complement 
assign qve = ~QVE;  //complement 
assign nbd = ~NBD;  //complement 
assign nbe = ~NBE;  //complement 
assign nbf = ~NBF;  //complement 
assign vab = ~VAB;  //complement 
assign TGB = ~tgb;  //complement 
assign wab = ~WAB;  //complement 
assign wbb = ~WBB;  //complement 
assign wcb = ~WCB;  //complement 
assign nba = ~NBA;  //complement 
assign nbb = ~NBB;  //complement 
assign nbc = ~NBC;  //complement 
assign nbg = ~NBG;  //complement 
assign nbh = ~NBH;  //complement 
assign nbi = ~NBI;  //complement 
assign nbj = ~NBJ;  //complement 
assign nbk = ~NBK;  //complement 
assign nbl = ~NBL;  //complement 
assign fba =  nba  ; 
assign FBA = ~fba;  //complement 
assign fbb =  nbb  ; 
assign FBB = ~fbb;  //complement 
assign fbc =  nbc  ; 
assign FBC = ~fbc;  //complement 
assign fbd =  nbd  ; 
assign FBD = ~fbd;  //complement 
assign fbe =  nbe  ; 
assign FBE = ~fbe;  //complement 
assign fbf =  nbf  ; 
assign FBF = ~fbf;  //complement 
assign wdb = ~WDB;  //complement 
assign web = ~WEB;  //complement 
assign wfb = ~WFB;  //complement 
assign fbg =  nbg  ; 
assign FBG = ~fbg;  //complement 
assign fbh =  nbh  ; 
assign FBH = ~fbh;  //complement 
assign fbi =  nbi  ; 
assign FBI = ~fbi;  //complement 
assign fbj =  nbj  ; 
assign FBJ = ~fbj;  //complement 
assign fbk =  nbk  ; 
assign FBK = ~fbk;  //complement 
assign fbl =  nbl  ; 
assign FBL = ~fbl;  //complement 
assign qvg = ~QVG;  //complement 
assign qvh = ~QVH;  //complement 
assign wgb = ~WGB;  //complement 
assign whb = ~WHB;  //complement 
assign saf = ~SAF;  //complement 
assign nkf = ~NKF;  //complement 
assign JPB =  QRD  ; 
assign jpb = ~JPB;  //complement 
assign jqb =  qau & qmc  ; 
assign JQB = ~jqb;  //complement 
assign JRB =  QAV  ; 
assign jrb = ~JRB;  //complement 
assign san = ~SAN;  //complement 
assign nkn = ~NKN;  //complement 
assign lbe = ~LBE;  //complement 
assign lbf = ~LBF;  //complement 
assign lbg = ~LBG;  //complement 
assign lbh = ~LBH;  //complement 
assign sav = ~SAV;  //complement 
assign raf = ~RAF;  //complement 
assign sce = ~SCE;  //complement 
assign scf = ~SCF;  //complement 
assign joe = ~JOE;  //complement 
assign jof = ~JOF;  //complement 
assign jog = ~JOG;  //complement 
assign joh = ~JOH;  //complement 
assign EAN =  AAN  ; 
assign ean = ~EAN;  //complement 
assign QJN =  QJO & sdm  ; 
assign qjn = ~QJN;  //complement 
assign scg = ~SCG;  //complement 
assign sch = ~SCH;  //complement 
assign QLF = ~qlf;  //complement 
assign QLG = ~qlg;  //complement 
assign QLL = ~qll;  //complement 
assign TBC =  QLE  ; 
assign tbc = ~TBC;  //complement 
assign kaf = ~KAF;  //complement 
assign okf = ~OKF;  //complement 
assign baf = ~BAF;  //complement 
assign ban = ~BAN;  //complement 
assign kan = ~KAN;  //complement 
assign kao = ~KAO;  //complement 
assign oif = ~OIF;  //complement 
assign oin = ~OIN;  //complement 
assign AAF = ~aaf;  //complement 
assign AAN = ~aan;  //complement 
assign ABF = ~abf;  //complement 
assign abn = ~ABN;  //complement 
assign tbo =  qlf  ; 
assign TBO = ~tbo;  //complement 
assign tbg =  qlf  ; 
assign TBG = ~tbg;  //complement 
assign tbi =  qlg  ; 
assign TBI = ~tbi;  //complement 
assign TBN =  QLE  ; 
assign tbn = ~TBN;  //complement 
assign TBM =  QLE  ; 
assign tbm = ~TBM;  //complement 
assign TBH =  QLI  ; 
assign tbh = ~TBH;  //complement 
assign ohf = ~OHF;  //complement 
assign ohn = ~OHN;  //complement 
assign okn = ~OKN;  //complement 
assign qfa = ~QFA;  //complement 
assign JBF =  AAW & aak & AAU  ; 
assign jbf = ~JBF;  //complement 
assign jdb =  qeb & qfb & qfc  ; 
assign JDB = ~jdb;  //complement 
assign lae = ~LAE;  //complement 
assign laf = ~LAF;  //complement 
assign lag = ~LAG;  //complement 
assign lah = ~LAH;  //complement 
assign ona = ~ONA;  //complement 
assign onb = ~ONB;  //complement 
assign daf = ~DAF;  //complement 
assign qfb = ~QFB;  //complement 
assign qfc = ~QFC;  //complement 
assign JKA =  QKC & qkb & qka  ; 
assign jka = ~JKA;  //complement 
assign JKB =  QKC & qkb & QKA  ; 
assign jkb = ~JKB;  //complement 
assign NLF =  RAF & QLJ & QKA  ; 
assign nlf = ~NLF;  //complement 
assign JKC =  QKC & QKB & qka  ; 
assign jkc = ~JKC;  //complement 
assign JKD =  QKC & QKB & QKA  ; 
assign jkd = ~JKD;  //complement 
assign qka = ~QKA;  //complement 
assign qkb = ~QKB;  //complement 
assign qkc = ~QKC;  //complement 
assign thi = ~THI;  //complement 
assign thj = ~THJ;  //complement 
assign thk = ~THK;  //complement 
assign thl = ~THL;  //complement 
assign ncd = ~NCD;  //complement 
assign nce = ~NCE;  //complement 
assign ncf = ~NCF;  //complement 
assign vac = ~VAC;  //complement 
assign TGC = ~tgc;  //complement 
assign wac = ~WAC;  //complement 
assign wbc = ~WBC;  //complement 
assign wcc = ~WCC;  //complement 
assign nca = ~NCA;  //complement 
assign ncb = ~NCB;  //complement 
assign ncc = ~NCC;  //complement 
assign ncg = ~NCG;  //complement 
assign nch = ~NCH;  //complement 
assign nci = ~NCI;  //complement 
assign ncj = ~NCJ;  //complement 
assign nck = ~NCK;  //complement 
assign ncl = ~NCL;  //complement 
assign fca =  nca  ; 
assign FCA = ~fca;  //complement 
assign fcb =  ncb  ; 
assign FCB = ~fcb;  //complement 
assign fcc =  ncc  ; 
assign FCC = ~fcc;  //complement 
assign fcd =  ncd  ; 
assign FCD = ~fcd;  //complement 
assign fce =  nce  ; 
assign FCE = ~fce;  //complement 
assign fcf =  ncf  ; 
assign FCF = ~fcf;  //complement 
assign qvf = ~QVF;  //complement 
assign fcg =  ncg  ; 
assign FCG = ~fcg;  //complement 
assign fch =  nch  ; 
assign FCH = ~fch;  //complement 
assign fci =  nci  ; 
assign FCI = ~fci;  //complement 
assign fcj =  ncj  ; 
assign FCJ = ~fcj;  //complement 
assign fck =  nck  ; 
assign FCK = ~fck;  //complement 
assign fcl =  ncl  ; 
assign FCL = ~fcl;  //complement 
assign wdc = ~WDC;  //complement 
assign wec = ~WEC;  //complement 
assign wfc = ~WFC;  //complement 
assign wgc = ~WGC;  //complement 
assign whc = ~WHC;  //complement 
assign qvi = ~QVI;  //complement 
assign qvj = ~QVJ;  //complement 
assign sag = ~SAG;  //complement 
assign nkg = ~NKG;  //complement 
assign JPC =  QRD  ; 
assign jpc = ~JPC;  //complement 
assign jqc =  qau & qmc  ; 
assign JQC = ~jqc;  //complement 
assign JRC =  QAV  ; 
assign jrc = ~JRC;  //complement 
assign sao = ~SAO;  //complement 
assign lbi = ~LBI;  //complement 
assign lbj = ~LBJ;  //complement 
assign lbk = ~LBK;  //complement 
assign lbl = ~LBL;  //complement 
assign saw = ~SAW;  //complement 
assign rag = ~RAG;  //complement 
assign sci = ~SCI;  //complement 
assign scj = ~SCJ;  //complement 
assign joi = ~JOI;  //complement 
assign joj = ~JOJ;  //complement 
assign jok = ~JOK;  //complement 
assign jol = ~JOL;  //complement 
assign qgb = ~QGB;  //complement 
assign sck = ~SCK;  //complement 
assign scl = ~SCL;  //complement 
assign kag = ~KAG;  //complement 
assign okg = ~OKG;  //complement 
assign bag = ~BAG;  //complement 
assign bao = ~BAO;  //complement 
assign EAO =  AAO  ; 
assign eao = ~EAO;  //complement 
assign oig = ~OIG;  //complement 
assign oio = ~OIO;  //complement 
assign AAG = ~aag;  //complement 
assign AAO = ~aao;  //complement 
assign ABG = ~abg;  //complement 
assign abo = ~ABO;  //complement 
assign qid = ~QID;  //complement 
assign qja = ~QJA;  //complement 
assign qjb = ~QJB;  //complement 
assign ohg = ~OHG;  //complement 
assign oho = ~OHO;  //complement 
assign oko = ~OKO;  //complement 
assign qga = ~QGA;  //complement 
assign JBG =  AAW & AAV & aaj  ; 
assign jbg = ~JBG;  //complement 
assign NLG =  RAG & QLJ  ; 
assign nlg = ~NLG;  //complement 
assign lai = ~LAI;  //complement 
assign laj = ~LAJ;  //complement 
assign lak = ~LAK;  //complement 
assign lal = ~LAL;  //complement 
assign qxd = ~QXD;  //complement 
assign qxe = ~QXE;  //complement 
assign qxf = ~QXF;  //complement 
assign ola = ~OLA;  //complement 
assign ooa = ~OOA;  //complement 
assign ndd = ~NDD;  //complement 
assign nde = ~NDE;  //complement 
assign ndf = ~NDF;  //complement 
assign vad = ~VAD;  //complement 
assign TGD = ~tgd;  //complement 
assign wad = ~WAD;  //complement 
assign wbd = ~WBD;  //complement 
assign wcd = ~WCD;  //complement 
assign nda = ~NDA;  //complement 
assign ndb = ~NDB;  //complement 
assign ndc = ~NDC;  //complement 
assign ndg = ~NDG;  //complement 
assign ndh = ~NDH;  //complement 
assign ndi = ~NDI;  //complement 
assign ndj = ~NDJ;  //complement 
assign ndk = ~NDK;  //complement 
assign ndl = ~NDL;  //complement 
assign fda =  nda  ; 
assign FDA = ~fda;  //complement 
assign fdb =  ndb  ; 
assign FDB = ~fdb;  //complement 
assign fdc =  ndc  ; 
assign FDC = ~fdc;  //complement 
assign fdd =  ndd  ; 
assign FDD = ~fdd;  //complement 
assign fde =  nde  ; 
assign FDE = ~fde;  //complement 
assign fdf =  ndf  ; 
assign FDF = ~fdf;  //complement 
assign fdg =  ndg  ; 
assign FDG = ~fdg;  //complement 
assign fdh =  ndh  ; 
assign FDH = ~fdh;  //complement 
assign fdi =  ndi  ; 
assign FDI = ~fdi;  //complement 
assign fdj =  ndj  ; 
assign FDJ = ~fdj;  //complement 
assign fdk =  ndk  ; 
assign FDK = ~fdk;  //complement 
assign fdl =  ndl  ; 
assign FDL = ~fdl;  //complement 
assign wdd = ~WDD;  //complement 
assign wed = ~WED;  //complement 
assign wfd = ~WFD;  //complement 
assign qwb = ~QWB;  //complement 
assign QYA =  QWA  |  QWB  |  QWC  |  QWD  ;
assign qya = ~QYA;  //complement 
assign wgd = ~WGD;  //complement 
assign whd = ~WHD;  //complement 
assign qwd = ~QWD;  //complement 
assign qvk = ~QVK;  //complement 
assign sah = ~SAH;  //complement 
assign nkh = ~NKH;  //complement 
assign qwf = ~QWF;  //complement 
assign sap = ~SAP;  //complement 
assign QJK =  QJF & sam  ; 
assign qjk = ~QJK;  //complement 
assign QJL =  QJF & sam  ; 
assign qjl = ~QJL;  //complement 
assign QJM =  QJF & sam  ; 
assign qjm = ~QJM;  //complement 
assign qmc = ~QMC;  //complement 
assign qhb = ~QHB;  //complement 
assign sax = ~SAX;  //complement 
assign rah = ~RAH;  //complement 
assign qwc = ~QWC;  //complement 
assign QJF = ~qjf;  //complement 
assign QJO = ~qjo;  //complement 
assign QJP = ~qjp;  //complement 
assign qlh = ~QLH;  //complement 
assign qle = ~QLE;  //complement 
assign qwa = ~QWA;  //complement 
assign qli = ~QLI;  //complement 
assign qlj = ~QLJ;  //complement 
assign qlk = ~QLK;  //complement 
assign QYB =  QWE  |  QWF  |  QWG  |  QWH  ;
assign qyb = ~QYB;  //complement 
assign qwe = ~QWE;  //complement 
assign qza = ~QZA;  //complement 
assign qzb = ~QZB;  //complement 
assign qzc = ~QZC;  //complement 
assign qzd = ~QZD;  //complement 
assign TBE =  QLI  ; 
assign tbe = ~TBE;  //complement 
assign qwg = ~QWG;  //complement 
assign qze = ~QZE;  //complement 
assign qzf = ~QZF;  //complement 
assign qzg = ~QZG;  //complement 
assign qzh = ~QZH;  //complement 
assign qwh = ~QWH;  //complement 
assign kah = ~KAH;  //complement 
assign kap = ~KAP;  //complement 
assign okh = ~OKH;  //complement 
assign bah = ~BAH;  //complement 
assign bap = ~BAP;  //complement 
assign oih = ~OIH;  //complement 
assign oip = ~OIP;  //complement 
assign AAH = ~aah;  //complement 
assign AAP = ~aap;  //complement 
assign ABH = ~abh;  //complement 
assign abp = ~ABP;  //complement 
assign ohh = ~OHH;  //complement 
assign ohp = ~OHP;  //complement 
assign okp = ~OKP;  //complement 
assign qha = ~QHA;  //complement 
assign JBH =  AAW & AAV & AAU  ; 
assign jbh = ~JBH;  //complement 
assign NLH =  RAH & QLJ  ; 
assign nlh = ~NLH;  //complement 
assign qug = ~QUG;  //complement 
assign quh = ~QUH;  //complement 
assign qui = ~QUI;  //complement 
assign olb = ~OLB;  //complement 
assign qxg = ~QXG;  //complement 
assign quj = ~QUJ;  //complement 
assign quk = ~QUK;  //complement 
assign qul = ~QUL;  //complement 
assign qum = ~QUM;  //complement 
assign qun = ~QUN;  //complement 
assign qxa = ~QXA;  //complement 
assign qxb = ~QXB;  //complement 
assign qxc = ~QXC;  //complement 
assign oja = ~OJA;  //complement 
assign ojb = ~OJB;  //complement 
assign ojc = ~OJC;  //complement 
assign ojd = ~OJD;  //complement 
assign qxh = ~QXH;  //complement 
assign oje = ~OJE;  //complement 
assign ojf = ~OJF;  //complement 
assign ojg = ~OJG;  //complement 
assign ojh = ~OJH;  //complement 
assign oji = ~OJI;  //complement 
assign ojj = ~OJJ;  //complement 
assign qmb = ~QMB;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign icq = ~ICQ; //complement 
assign icr = ~ICR; //complement 
assign ics = ~ICS; //complement 
assign ict = ~ICT; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign iga = ~IGA; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign iic = ~IIC; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign iki = ~IKI; //complement 
assign ikj = ~IKJ; //complement 
assign ikk = ~IKK; //complement 
assign ikl = ~IKL; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ild = ~ILD; //complement 
assign ile = ~ILE; //complement 
assign ilf = ~ILF; //complement 
assign ilg = ~ILG; //complement 
assign ilh = ~ILH; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign imh = ~IMH; //complement 
assign ixa = ~IXA; //complement 
always@(posedge IZZ )
   begin 
 SAA <=  SAA & tca & qid  |  AAA & TCA  |  DAA & QID  ; 
 NKA <=  NKA & SDM & qhe  |  NJM & QJL  |  AAA & QHE  ; 
 SAI <=  SAI & tca  |  AAI & TCB  ; 
 NKI <=  NKI & SDM & qhe  |  NJG & QJN  |  AAI & QHE  ; 
 QAU <= QAH ; 
 QAV <= QAH ; 
 SAQ <=  SAQ & tcc  |  ABA & TCC  ; 
 RAA <=  RAA & SFM & qhg  |  QZA & QJK  |  ABA & QHG  ; 
 QLA <=  SAJ & SAP  |  SAK & SAQ  |  SAL & SAR  ; 
 QLB <=  SAM & SAS  |  SAN & SAT  |  SBB & SBC  ; 
 QAD <= QAC ; 
 QAE <= QAD ; 
 QAF <= QAE ; 
 QAG <= QAF ; 
 QAH <= QAG ; 
 QAI <= QAH ; 
 QAJ <= QAI ; 
 QAK <= QAJ ; 
 QAL <= QAK ; 
 QAM <= QAL ; 
 QAN <= QAM ; 
 QAO <= QAN ; 
 QAP <= QAO ; 
 QAQ <= QAP ; 
 SBA <=  SBA & tcd  |  ABI & TCD  ; 
 OMF <=  SBA & tcd  |  ABI & TCD  ; 
 KAA <=  IAA & TBA  |  SAA & TBB  |  SAQ & TBC  |  NKA & TBD  |  NLA  ; 
 KAI <=  IAI & TBA  |  SAI & TBB  |  SBA & TBM  |  NKI & TBD  ; 
 OKA <=  ICA & TAA  |  IBA & TAB  |  KAA & TAC  |  BAA & TAD  |  JOA  ; 
 BAA <=  AAA & TDA  |  BAA & tda  ; 
 BAI <=  AAI & TDA  |  BAI & tda  ; 
 OIA <=  ABA & tib  |  IBA & TIB  ; 
 OII <=  ABI & tib  |  IBI & TIB  ; 
 aaa <= ica ; 
 aai <= ici ; 
 aba <= aaa ; 
 abi <= aai ; 
 qia <=  qla & qlb  |  aaq  |  qib  ; 
 qie <=  qla & qlb  |  aaq  |  qib  ; 
 DAA <= IDA ; 
 ojk <= qma ; 
 ojl <= qma ; 
 AAT <= ICA ; 
 OHA <=  AAA & tia  |  IAA & TIA  ; 
 OHI <=  AAI & tia  |  IAI & TIA  ; 
 OKI <=  ICI & TAI  |  IBI & TAF  |  KAI & TAG  |  BAI & TAH  |  JOI  ; 
 QAA <=  JAA & JBA  ; 
 OKQ <= ICQ ; 
 qic <= ieg ; 
 QMA <= IGA ; 
 OLC <= SAI ; 
 QAB <=  QAB & aas & jma  |  QAA  ; 
 QOB <=  QOB & qod & jmb  |  QOA  ; 
 QOF <=  QOB & qod & jmb  |  QOA  ; 
 OMB <=  QAE  |  QGB  |  QCA  ; 
 aaq <= icq ; 
 abq <= aaq ; 
 OMC <= QAM ; 
 OMD <= QAQ ; 
 QAC <=  QAB & AAS  ; 
 QAS <=  QAR & qib  ; 
 QAR <=  QAR & QIB & jmb  |  QAQ  ; 
 QIB <=  IEC & qic & qqb  ; 
 had <=  jna  ; 
 hag <=  jnb  |  jnd  ; 
 haj <=  jnc  |  jne  |  jnf  ; 
 SAB <=  SAB & tca & qid  |  AAB & TCA  |  DAB & QID  ; 
 NKB <=  NKB & SDM & qhe  |  NJN & QJL  |  AAB & QHE  ; 
 SAJ <=  SAJ & tcb  |  AAJ & TCB  |  QJC  ; 
 NKJ <=  NKJ & SEM & qhe  |  NJH & QJN  |  AAJ & QHE  ; 
 SAR <=  SAR & tcc  |  ABB & TCC  ; 
 RAB <=  RAB & SFM & qhg  |  QZB & QJK  |  ABB & QHG  ; 
 QLC <=  QBC  |  QEA  ; 
 QLD <=  JDA  |  JDB  ; 
 QBB <= QBA ; 
 QBC <= QBB ; 
 QBD <= QBC ; 
 QBE <= QBD ; 
 QBF <= QBE ; 
 QBG <= QBF ; 
 QBH <= QBG ; 
 QBI <= QBH ; 
 KAB <=  IAB & TBA  |  SAB & TBB  |  SAR & TBC  |  NKB & TBD  |  NLB  ; 
 KAJ <=  IAJ & TBA  |  SAJ & TBB  |  SBB & TBM  |  NKJ & TBD  ; 
 OKB <=  ICB & TAA  |  IBB & TAB  |  KAB & TAC  |  BAB & TAD  |  JOB  ; 
 BAB <=  AAB & TDA  |  BAB & tda  ; 
 BAJ <=  AAJ & TDA  |  BAJ & tda  ; 
 OIB <=  ABB & tib  |  IBB & TIB  ; 
 OIJ <=  ABJ & tib  |  IBJ & TIB  ; 
 aab <= icb ; 
 aaj <= icj ; 
 abb <= aab ; 
 AAU <= ICJ ; 
 DAB <= IDB ; 
 QJE <= IFD ; 
 qoa <= jaa ; 
 ACJ <= ICJ ; 
 OHB <=  AAB & tia  |  IAB & TIA  ; 
 OHJ <=  ACJ & tia  |  IAJ & TIA  ; 
 OKJ <=  ICJ & TAI  |  IBJ & TAF  |  KAJ & TAG  |  BAJ & TAH  |  JOJ  ; 
 QBA <=  JAA & JBB  ; 
 OKR <=  ICR  ; 
 SBB <=  SBB & tcd  |  ABJ & TCD  |  IEE  ; 
 QBJ <=  QBJ & aas & jmb  |  QBI  ; 
 QJC <=  IFA  |  IFB  ; 
 aar <= icr ; 
 abr <= aar ; 
 abj <= aaj ; 
 QBK <=  QBJ & AAS  ; 
 QTB <=  QSB  |  QSD  ; 
 QUC <= QUB ; 
 QUD <= QUC ; 
 QUE <= QUD ; 
 QUF <= QUE ; 
 QUA <=  QSA  |  QSC  ; 
 QUB <=  QUA  ; 
 qsa <=  qra  |  QQB  |  QQC  ; 
 qsb <=  qra  |  qqb  |  QQC  ; 
 qsc <=  qrc  |  QQB  ; 
 qsd <=  qrc  |  qqb  ; 
 hab <=  nba  ; 
 hae <=  jna  |  nbd  ; 
 hah <=  jnb  |  jnd  |  nbg  ; 
 hak <=  jnc  |  jne  |  jnf  |  nbj  ; 
 SAC <=  SAC & tca & qid  |  AAC & TCA  |  DAC & QID  ; 
 NKC <=  NKC & SDM & qhe  |  NJA & QJL  |  AAC & QHE  ; 
 QPA <= QRA ; 
 QPB <= QSE ; 
 SAK <=  SAK & tcb  |  AAK & TCB  |  QJD & QJJ  ; 
 NKK <=  NKK & SEM & qhe  |  NJI & QJN  |  AAK & QHE  ; 
 QRA <= QQA ; 
 QRB <= QQB ; 
 QRC <= QQC ; 
 QSE <= QRC ; 
 SAS <=  SAS & tcc  |  ABC & TCC  ; 
 RAC <=  RAC & SFM & qhg  |  QZC & QJK  |  ABC & QHG  ; 
 TEA <= QRA ; 
 TEB <= QRA ; 
 TEC <= QRA ; 
 TED <= QRA ; 
 QRD <=  QQB & QRA  |  QQB & QRE  ; 
 QRE <=  QQC & QRA  ; 
 QHC <= aba & QHB ; 
 QHD <= aba & QHB ; 
 QAT <= QAI ; 
 QHE <= ABA & QHB ; 
 QHF <= ABA & QHB ; 
 QHG <= ABA & QHB ; 
 QHH <= ABA & QHB ; 
 KAC <=  IAC & TBA  |  SAC & TBB  |  SAS & TBC  |  NKC & TBD  |  NLC  ; 
 KAK <=  IAK & TBA  |  SAK & TBB  |  SBC & TBM  |  NKK & TBD  ; 
 OKC <=  ICC & TAA  |  IBC & TAB  |  KAC & TAC  |  BAC & TAD  |  JOC  ; 
 BAC <=  AAC & TDA  |  BAC & tda  ; 
 BAK <=  AAK & TDA  |  BAK & tda  ; 
 TIA <= QCA ; 
 TIB <= QCA ; 
 OIC <=  ABC & tib  |  IBC & TIB  ; 
 OIK <=  ABK & tib  |  IBK & TIB  ; 
 aac <= icc ; 
 aak <= ick ; 
 abc <= aac ; 
 AAV <= ICK ; 
 SBC <=  SBC & tcd  |  ABK & TCD  ; 
 DAC <= IDC ; 
 QJD <= IFC ; 
 ACK <= ICK ; 
 abk <= aak ; 
 OHC <=  AAC & tia  |  IAC & TIA  ; 
 OHK <=  ACK & tia  |  IAK & TIA  ; 
 OKK <=  ICK & TAE  |  IBK & TAF  |  KAK & TAG  |  BAK & TAH  |  JOK  ; 
 QCA <=  JAA & JBC  ; 
 QJG <= IEF ; 
 QJH <= QJG ; 
 QJI <= QJH ; 
 QJJ <= QJI ; 
 OKS <=  ICS & qbj & qab  |  QBA  |  QAS  ; 
 QCB <=  QCB & QIB & jma  |  QCA  ; 
 aas <= ics ; 
 QQA <= IIA ; 
 QQB <= IIB ; 
 QQC <= IIC ; 
 QCC <=  QCB & qib  ; 
 abs <= aas ; 
 OME <=  QCA  |  QAQ  ; 
 TFA <= QTB & PAA ; 
 TFB <= QTB & PAB ; 
 TFC <= QTB & PAC ; 
 TFD <= QTB & PAD ; 
 hac <=  nba  |  nbb  ; 
 haf <=  jna  |  nbd  |  nbe  ; 
 hai <=  jnb  |  jnd  |  nbg  |  nbh  ; 
 hal <=  jnc  |  jne  |  jnf  |  nbj  |  nbk  ; 
 PAA <=  PAA & qpa & qpb  |  LBM & QPA  |  PAD & QPB  ; 
 PAB <=  PAB & qpa & qpb  |  LBN & QPA  |  PAA & QPB  ; 
 PAC <=  PAC & qpa & qpb  |  LBO & QPA  |  PAB & QPB  ; 
 PAD <=  PAD & qpa & qpb  |  LBP & QPA  |  PAC & QPB  ; 
 pba <= paa ; 
 pca <= pba ; 
 pbb <= pab ; 
 pcb <= pbb ; 
 pbc <= pac ; 
 pcc <= pbc ; 
 pbd <= pad ; 
 pcd <= pbd ; 
 SAD <=  SAD & tca & qid  |  AAD & TCA  |  DAD & QID  ; 
 NKD <=  NKD & SDM & qhe  |  NJB & QJL  |  AAD & QHE  ; 
 SAL <=  SAL & tcb  |  AAL & TCB  |  QJE  ; 
 NKL <=  NKL & SEM & qhe  |  NJJ & QJN  |  AAL & QHE  ; 
 SAT <=  SAT & tcc  |  ABD & TCC  ; 
 RAD <=  RAD & SFM & qhg  |  QZD & QJM  |  ABD & QHG  ; 
 QNA <=  QSE & PAD & qpb  |  QPB & PAC  ; 
 QNB <=  QSE & PAD & qpb  |  QPB & PAC  ; 
 QNC <=  QSE & PAD & qpb  |  QPB & PAC  ; 
 LBM <= LAM ; 
 LBN <= LAN ; 
 LBO <= LAO ; 
 LBP <= LAP ; 
 QDD <= QDC ; 
 tbb <= tbc ; 
 KAL <=  IAL & TBP  |  SAL & TBO  |  NKL & TBQ  ; 
 KAM <=  IAM & TBP  |  SAM & TBO  |  NKM & TBQ  ; 
 OKD <=  ICD & TAA  |  IBD & TAB  |  KAD & TAC  |  BAD & TAD  |  JOD  ; 
 BAD <=  AAD & TDA  |  BAD & tda  ; 
 BAL <=  AAL & TDA  |  BAL & tda  ; 
 KAD <=  IAD & TBA  |  SAD & TBB  |  SAT & TBC  |  NKD & TBD  |  NLD  ; 
 OID <=  ABD & tib  |  IBD & TIB  ; 
 OIL <=  ABL & tib  |  IBL & TIB  ; 
 aad <= icd ; 
 aal <= icl ; 
 abd <= aad ; 
 AAW <= ICL ; 
 DAD <= IDD ; 
 QOD <= QOC ; 
 ACL <= ICL ; 
 abl <= aal ; 
 OHD <=  AAD & tia  |  IAD & TIA  ; 
 OHL <=  ACL & tia  |  IAL & TIA  ; 
 OKL <=  ICL & TAE  |  IBL & TAF  |  KAL & TAG  |  BAL & TAH  |  JOL  ; 
 QDA <=  JAA & JBD  ; 
 OKT <=  ICT  |  JCF  |  JCG  ; 
 QOC <=  ICT  |  JCF  |  JCG  ; 
 QDB <=  QDB & qib & jma  |  QDA  ; 
 OMA <=  QDA  |  JGA  ; 
 QDC <=  QDB & QIB  ; 
 LAM <= IJA ; 
 LAN <= IJB ; 
 LAO <= IJC ; 
 LAP <= IJD ; 
 THA <= QUC & PCA ; 
 THB <= QUC & PCB ; 
 THC <= QUC & PCC ; 
 THD <= QUC & PCD ; 
 QVD <=  MAA & THA  |  MAB & THB  |  MAC & THC  |  MAD & THD  ; 
 THE <= QUC & PCA ; 
 THF <= QUC & PCB ; 
 THG <= QUC & PCC ; 
 THH <= QUC & PCD ; 
 NAD <= GAD & tea |  LBD & TEA ; 
 NAE <= GAE & tea |  LBE & TEA ; 
 NAF <= GAF & tea |  LBF & TEA ; 
 VAA <=  TFA  |  TGA  ; 
 tga <=  tfa  ; 
 WAA <= WAA & tfa |  QXA & TFA ; 
 WBA <= WBA & tfa |  QXB & TFA ; 
 WCA <= WCA & tfa |  QXC & TFA ; 
 NAA <= GAA & tea |  LBA & TEA ; 
 NAB <= GAB & tea |  LBB & TEA ; 
 NAC <= GAC & tea |  LBC & TEA ; 
 NAG <= GAG & tea |  LBG & TEA ; 
 NAH <= GAH & tea |  LBH & TEA ; 
 NAI <= GAI & tea |  LBI & TEA ; 
 NAJ <= GAJ & tea |  LBJ & TEA ; 
 NAK <= GAK & tea |  LBK & TEA ; 
 NAL <= GAL & tea |  LBL & TEA ; 
 WDA <= WDA & tfa |  QXD & TFA ; 
 WEA <= WEA & tfa |  QXE & TFA ; 
 WFA <= WFA & tfa |  QXF & TFA ; 
 WGA <= WGA & tfa |  QXG & TFA ; 
 WHA <= WHA & tfa |  QXH & TFA ; 
 NEA <= NAA ; 
 NEB <= NAB ; 
 NEC <= NAC ; 
 NED <= NAD ; 
 NEE <= NAE ; 
 NEF <= NAF ; 
 NEG <= NAG ; 
 NEH <= NAH ; 
 NEI <= NAI ; 
 NEJ <= NAJ ; 
 NEK <= NAK ; 
 NEL <= NAL ; 
 NFA <= NEA ; 
 NFB <= NEB ; 
 NFC <= NEC ; 
 NFD <= NED ; 
 NHM <=  THB  |  THD  ; 
 NHN <=  THD  |  THC  ; 
 SAE <=  SAE & tce & qid  |  AAE & TCE  |  DAE & QID  ; 
 NKE <=  NKE & SDM & qhf  |  NJC & QJL  |  AAE & QHF  ; 
 SAM <=  SAM & tce  |  EAM & TCE  |  QJP  ; 
 SDM <=  SAM & tce  |  EAM & TCE  |  QJP  ; 
 SEM <=  SAM & tce  |  EAM & TCE  |  QJP  ; 
 NKM <=  NKM & SEM & qhf  |  NJK & QJN  |  AAM & QHF  ; 
 LBA <= LAA ; 
 LBB <= LAB ; 
 LBC <= LAC ; 
 LBD <= LAD ; 
 SAU <=  QIB  ; 
 RAE <=  RAE & SFM & qhh  |  QZE & QJM  |  ABE & QHH  ; 
 SCA <=  SCA & jqa  |  LBA & JPA  |  ABA & JRA  ; 
 SCB <=  SCB & jqa  |  LBB & JPA  |  ABB & JRA  ; 
 JOA <= QBF & SCA ; 
 JOB <= QBF & SCB ; 
 JOC <= QBF & SCC ; 
 JOD <= QBF & SCD ; 
 QEB <= QEA ; 
 SCC <=  SCC & jqa  |  LBC & JPA  |  ABC & JRA  ; 
 SCD <=  SCD & jqa  |  LBD & JPA  |  ABD & JRA  ; 
 NHE <= NGE ; 
 NHF <= NGF ; 
 NHG <= NGG ; 
 NHH <= NGH ; 
 NIA <= NHA ; 
 NIB <= NHB ; 
 NIC <= NHC ; 
 NID <= NHD ; 
 NGA <= NFA ; 
 NGB <= NFB ; 
 NGC <= NFC ; 
 NGD <= NFD ; 
 NGE <= NFE ; 
 NGF <= NFF ; 
 NGG <= NFG ; 
 NGH <= NFH ; 
 NIE <= NHE ; 
 NIF <= NHF ; 
 NIG <= NHG ; 
 NIH <= NHH ; 
 NFI <= NEI ; 
 NFJ <= NEJ ; 
 NFK <= NEK ; 
 NFL <= NEL ; 
 NGI <= NFI ; 
 NGJ <= NFJ ; 
 NGK <= NFK ; 
 NGL <= NFL ; 
 NII <= NHI ; 
 NIJ <= NHJ ; 
 NIK <= NHK ; 
 NIL <= NHL ; 
 NFE <= NEE ; 
 NFF <= NEF ; 
 NFG <= NEG ; 
 NFH <= NEH ; 
 NHI <= NGI ; 
 NHJ <= NGJ ; 
 NHK <= NGK ; 
 NHL <= NGL ; 
 KAE <=  IAE & TBP  |  SAE & TBO  |  SAU & TBN  |  NKE & TBI  |  NLE  ; 
 OKE <=  ICE & TAJ  |  IBE & TAB  |  KAE & TAC  |  BAE & TAD  |  JOE  ; 
 BAE <=  AAE & TDA  |  BAE & tda  ; 
 BAM <=  EAM & TDA  |  BAM & tda  ; 
 SFM <=  SFM & tce  |  EAM & TCE  |  QJP  ; 
 OIE <=  ABE & tib  |  IBE & TIB  ; 
 OIM <=  ABM & tib  |  IBM & TIB  ; 
 aae <= ice ; 
 aam <= icm ; 
 abe <= aae ; 
 AAX <= ICM ; 
 NHA <= NGA ; 
 NHB <= NGB ; 
 NHC <= NGC ; 
 NHD <= NGD ; 
 DAE <= IDE ; 
 abm <= aam ; 
 OHE <=  AAE & tia  |  IAE & TIA  ; 
 OHM <=  AAM & tia  |  IAM & TIA  ; 
 OKM <=  ICM & TAE  |  IBM & TAF  |  KAM & TAG  |  BAM & TAH  ; 
 QEA <=  JAA & JBE  ; 
 LAA <= IKA ; 
 LAB <= IKB ; 
 LAC <= IKC ; 
 LAD <= IKD ; 
 NJA <= NIA ; 
 NJB <= NIB ; 
 NJC <= NIC ; 
 NJD <= NID ; 
 NJE <= NIE ; 
 NJF <= NIF ; 
 NJG <= NIG ; 
 NJH <= NIH ; 
 NJI <= NII ; 
 NJJ <= NIJ ; 
 NJK <= NIK ; 
 NJL <= NIL ; 
 NIM <= NHM ; 
 NIN <= NHN ; 
 NJM <= NIM ; 
 NJN <= NIN ; 
 QVE <=  MBA & THA  |  MBB & THB  |  MBC & THC  |  MBD & THD  ; 
 NBD <= FAM & teb |  LBD & TEB ; 
 NBE <= FAN & teb |  LBE & TEB ; 
 NBF <= FAF & teb |  LBF & TEB ; 
 VAB <=  TFB  |  TGB  ; 
 tgb <=  tfb  ; 
 WAB <= WAB & tfb |  QXA & TFB ; 
 WBB <= WBB & tfb |  QXB & TFB ; 
 WCB <= WCB & tfb |  QXC & TFB ; 
 NBA <= FAA & teb |  LBA & TEB ; 
 NBB <= FAB & teb |  LBB & TEB ; 
 NBC <= FAC & teb |  LBC & TEB ; 
 NBG <= FAG & teb |  LBG & TEB ; 
 NBH <= FAH & teb |  LBH & TEB ; 
 NBI <= FAI & teb |  LBI & TEB ; 
 NBJ <= FAJ & teb |  LBJ & TEB ; 
 NBK <= FAK & teb |  LBK & TEB ; 
 NBL <= FAL & teb |  LBL & TEB ; 
 WDB <= WDB & tfb |  QXD & TFB ; 
 WEB <= WEB & tfb |  QXE & TFB ; 
 WFB <= WFB & tfb |  QXF & TFB ; 
 QVG <=  MDA & THE  |  MDB & THF  |  MDC & THG  |  MDD & THH  ; 
 QVH <=  MEA & THE  |  MEB & THF  |  MEC & THG  |  MED & THH  ; 
 WGB <= WGB & tfb |  QXG & TFB ; 
 WHB <= WHB & tfb |  QXH & TFB ; 
 SAF <=  SAF & tce & qid  |  AAF & TCE  |  DAF & QID  ; 
 NKF <=  NKF & SDM & qhf  |  NJD & QJL  |  AAF & QHF  ; 
 SAN <=  SAN & tcb  |  EAN & TCB  |  QID  ; 
 NKN <=  NKN & SEM & qhf  |  NJL & QJN  |  AAN & QHF  ; 
 LBE <= LAE ; 
 LBF <= LAF ; 
 LBG <= LAG ; 
 LBH <= LAH ; 
 SAV <=  SAV & tcc & jkc  |  ABF & TCC  |  JKD  ; 
 RAF <=  RAF & SFM & qhh  |  QZF & QJM  |  ABF & QHH  ; 
 SCE <=  SCE & jqb  |  LBE & JPB  |  ABE & JRB  ; 
 SCF <=  SCF & jqb  |  LBF & JPB  |  ABF & JRB  ; 
 JOE <= QBF & SCE ; 
 JOF <= QBF & SCF ; 
 JOG <= QBF & SCG ; 
 JOH <= QBF & SCH ; 
 SCG <=  SCG & jqb  |  LBG & JPB  |  ABG & JRB  ; 
 SCH <=  SCH & jqb  |  LBH & JPB  |  ABH & JRB  ; 
 qlf <= tbc ; 
 qlg <= tbe ; 
 qll <= tbe ; 
 KAF <=  IAF & TBF  |  SAF & TBG  |  SAV & TBH  |  NKF & TBI  |  NLF  ; 
 OKF <=  ICF & TAJ  |  IBF & TAB  |  KAF & TAC  |  BAF & TAD  |  JOF  ; 
 BAF <=  AAF & TDA  |  BAF & tda  ; 
 BAN <=  EAN & TDA  |  BAN & tda  ; 
 KAN <=  IAN & TBF  |  SAN & TBG  |  NKN & TBQ  ; 
 KAO <=  IAO & TBF  |  SAO & TBG  ; 
 OIF <=  ABF & tib  |  IBF & TIB  ; 
 OIN <=  ABN & tib  |  IBN & TIB  ; 
 aaf <= icf ; 
 aan <= icn ; 
 abf <= aaf ; 
 ABN <= AAN ; 
 OHF <=  AAF & tia  |  IAF & TIA  ; 
 OHN <=  AAN & tia  |  IAN & TIA  ; 
 OKN <=  ICN & TAE  |  IBN & TAF  |  KAN & TAG  |  BAN & TAH  ; 
 QFA <= JBF & JAA ; 
 LAE <= IKE ; 
 LAF <= IKF ; 
 LAG <= IKG ; 
 LAH <= IKH ; 
 ONA <= SAV ; 
 ONB <= SAV ; 
 DAF <= IDF ; 
 QFB <= QFA ; 
 QFC <= QFB ; 
 QKA <= IHA ; 
 QKB <= IHB ; 
 QKC <= IHC ; 
 THI <= QUC & PCA ; 
 THJ <= QUC & PCB ; 
 THK <= QUC & PCC ; 
 THL <= QUC & PCD ; 
 NCD <= FBD & tec |  LBD & TEC ; 
 NCE <= FBE & tec |  LBE & TEC ; 
 NCF <= FBF & tec |  LBF & TEC ; 
 VAC <=  TFC  |  TGC  ; 
 tgc <=  tfc  ; 
 WAC <= WAC & tfc |  QXA & TFC ; 
 WBC <= WBC & tfc |  QXB & TFC ; 
 WCC <= WCC & tfc |  QXC & TFC ; 
 NCA <= FBA & tec |  LBA & TEC ; 
 NCB <= FBB & tec |  LBB & TEC ; 
 NCC <= FBC & tec |  LBC & TEC ; 
 NCG <= FBG & tec |  LBG & TEC ; 
 NCH <= FBH & tec |  LBH & TEC ; 
 NCI <= FBI & tec |  LBI & TEC ; 
 NCJ <= FBJ & tec |  LBJ & TEC ; 
 NCK <= FBK & tec |  LBK & TEC ; 
 NCL <= FBL & tec |  LBL & TEC ; 
 QVF <=  MCA & THE  |  MCB & THF  |  MCC & THG  |  MCD & THH  ; 
 WDC <= WDC & tfc |  QXD & TFC ; 
 WEC <= WEC & tfc |  QXE & TFC ; 
 WFC <= WFC & tfc |  QXF & TFC ; 
 WGC <= WGC & tfc |  QXG & TFC ; 
 WHC <= WHC & tfc |  QXH & TFC ; 
 QVI <=  MFA & THI  |  MFB & THJ  |  MFC & THK  |  MFD & THL  ; 
 QVJ <=  MGA & THI  |  MGB & THJ  |  MGC & THK  |  MGD & THL  ; 
 SAG <=  SAG & tca  |  AAG & TCA  ; 
 NKG <=  NKG & SDM & qhf  |  NJE & QJL  |  AAG & QHF  ; 
 SAO <=  SAO & tcb & qjb  |  EAO & TCB  |  QJA  ; 
 LBI <= LAI ; 
 LBJ <= LAJ ; 
 LBK <= LAK ; 
 LBL <= LAL ; 
 SAW <=  SAW & tcc & jka  |  ABG & TCC  |  JKB  ; 
 RAG <=  RAG & SFM & qhh  |  QZG & QJM  |  ABG & QHH  ; 
 SCI <=  SCI & jqc  |  LBI & JPC  |  ABI & JRC  ; 
 SCJ <=  SCJ & jqc  |  LBJ & JPC  |  ABJ & JRC  ; 
 JOI <= QBF & SCI ; 
 JOJ <= QBF & SCJ ; 
 JOK <= QBF & SCK ; 
 JOL <= QBF & SCL ; 
 QGB <= QGA ; 
 SCK <=  SCK & jqc  |  LBK & JPC  |  ABK & JRC  ; 
 SCL <=  SCL & jqc  |  LBL & JPC  |  ABL & JRC  ; 
 KAG <=  IAG & TBF  |  SAG & TBG  |  SAW & TBH  |  NKG & TBI  |  NLG  ; 
 OKG <=  ICG & TAJ  |  IBG & TAB  |  KAG & TAC  |  BAG & TAD  |  JOG  ; 
 BAG <=  AAG & TDA  |  BAG & tda  ; 
 BAO <=  EAO & TDA  |  BAO & tda  ; 
 OIG <=  ABG & tib  |  IBG & TIB  ; 
 OIO <=  ABO & tib  |  IBO & TIB  ; 
 aag <= icg ; 
 aao <= ico ; 
 abg <= aag ; 
 ABO <= AAO ; 
 QID <= IED ; 
 QJA <= IEA ; 
 QJB <= IEB ; 
 OHG <=  AAG & tia  |  IAG & TIA  ; 
 OHO <=  AAO & tia  |  IAO & TIA  ; 
 OKO <=  ICO & TAE  |  IBO & TAF  |  KAO & TAG  |  BAO & TAH  ; 
 QGA <=  JAA & JBG  ; 
 LAI <= IKI ; 
 LAJ <= IKJ ; 
 LAK <= IKK ; 
 LAL <= IKL ; 
 QXD <= ILD ; 
 QXE <= ILE ; 
 QXF <= ILF ; 
 OLA <= SAG ; 
 OOA <= SAW ; 
 NDD <= FCD & ted |  LBD & TED ; 
 NDE <= FCE & ted |  LBE & TED ; 
 NDF <= FCF & ted |  LBF & TED ; 
 VAD <=  TFD  |  TGD  ; 
 tgd <=  tfd  ; 
 WAD <= WAD & tfd |  QXA & TFD ; 
 WBD <= WBD & tfd |  QXB & TFD ; 
 WCD <= WCD & tfd |  QXC & TFD ; 
 NDA <= FCA & ted |  LBA & TED ; 
 NDB <= FCB & ted |  LBB & TED ; 
 NDC <= FCC & ted |  LBC & TED ; 
 NDG <= FCG & ted |  LBG & TED ; 
 NDH <= FCH & ted |  LBH & TED ; 
 NDI <= FCI & ted |  LBI & TED ; 
 NDJ <= FCJ & ted |  LBJ & TED ; 
 NDK <= FCK & ted |  LBK & TED ; 
 NDL <= FCL & ted |  LBL & TED ; 
 WDD <= WDD & tfd |  QXD & TFD ; 
 WED <= WED & tfd |  QXE & TFD ; 
 WFD <= WFD & tfd |  QXF & TFD ; 
 QWB <=  QUH & qve  |  quh & QVE  ; 
 WGD <= WGD & tfd |  QXG & TFD ; 
 WHD <= WHD & tfd |  QXH & TFD ; 
 QWD <=  QUJ & qvg  |  quj & QVG  ; 
 QVK <=  MHA & THI  |  MHB & THJ  |  MHC & THK  |  MHD & THL  ; 
 SAH <=  SAH & tca  |  AAH & TCA  ; 
 NKH <=  NKH & SDM & qhf  |  NJF & QJL  |  AAH & QHF  ; 
 QWF <=  QUL & qvi  |  qul & QVI  ; 
 SAP <=  SAP & tcb  |  AAP & TCB  ; 
 QMC <= QMB ; 
 QHB <= QHA ; 
 SAX <=  SAX & tcc  |  ABH & TCC  ; 
 RAH <=  RAH & SFM & qhh  |  QZH & QJM  |  ABH & QHH  ; 
 QWC <=  QUI & qvf  |  qui & QVF  ; 
 qjf <=  qya & qyb  |  quf  ; 
 qjo <=  qya & qyb  |  quf  ; 
 qjp <=  qya & qyb  |  quf  ; 
 QLH <=  QBF  |  aat & QFA  ; 
 QLE <=  QBF  |  aat & QFA  ; 
 QWA <=  QUG & qvd  |  qug & QVD  ; 
 QLI <= QFA & AAT ; 
 QLJ <= QFA & AAT ; 
 QLK <= QFA & AAT ; 
 QWE <=  QUK & qvh  |  quk & QVH  ; 
 QZA <= QWA ; 
 QZB <= QWB ; 
 QZC <= QWC ; 
 QZD <= QWD ; 
 QWG <=  QUM & qvj  |  qum & QVJ  ; 
 QZE <= QWE ; 
 QZF <= QWF ; 
 QZG <= QWG ; 
 QZH <= QWH ; 
 QWH <=  QUN & qvk  |  qun & QVK  ; 
 KAH <=  IAH & TBF  |  SAH & TBG  |  SAX & TBH  |  NKH & TBI  |  NLH  ; 
 KAP <=  IAP & TBF  |  SAP & TBG  ; 
 OKH <=  ICH & TAJ  |  IBH & TAB  |  KAH & TAC  |  BAH & TAD  |  JOH  ; 
 BAH <=  AAH & TDA  |  BAH & tda  ; 
 BAP <=  AAP & TDA  |  BAP & tda  ; 
 OIH <=  ABH & tib  |  IBH & TIB  ; 
 OIP <=  ABP & tib  |  IBP & TIB  ; 
 aah <= ich ; 
 aap <= icp ; 
 abh <= aah ; 
 ABP <= AAP ; 
 OHH <=  AAH & tia  |  IAH & TIA  ; 
 OHP <=  AAP & tia  |  IAP & TIA  ; 
 OKP <=  ICP & TAE  |  IBP & TAF  |  KAP & TAG  |  BAP & TAH  ; 
 QHA <=  JAA & JBH  ; 
 QUG <= IMA ; 
 QUH <= IMB ; 
 QUI <= IMC ; 
 OLB <= SAH ; 
 QXG <= ILG ; 
 QUJ <= IMD ; 
 QUK <= IME ; 
 QUL <= IMF ; 
 QUM <= IMG ; 
 QUN <= IMH ; 
 QXA <= ILA ; 
 QXB <= ILB ; 
 QXC <= ILC ; 
 OJA <= QMA ; 
 OJB <= QMA ; 
 OJC <= QMA ; 
 OJD <= QMA ; 
 QXH <= ILH ; 
 OJE <= QMA ; 
 OJF <= QMA ; 
 OJG <= QMA ; 
 OJH <= QMA ; 
 OJI <=  QMA  |  QAB  ; 
 OJJ <=  QMA  |  QAB  ; 
 QMB <=  QMA  |  QAB  ; 
 end 
end module
