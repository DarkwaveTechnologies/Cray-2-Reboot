module ar( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFF, 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 IHM, 
 IHN, 
 IHO, 
 IHP, 
 IIA, 
 IIB, 
 IIC, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IJF, 
 IKA, 
 IKB, 
 ILA, 
 IMA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OIJ, 
 OKA, 
 OKB, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 OMG, 
OMH ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFF; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 input IHM; 
 input IHN; 
 input IHO; 
 input IHP; 
 input IIA; 
 input IIB; 
 input IIC; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IJF; 
 input IKA; 
 input IKB; 
 input ILA; 
 input IMA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OIJ; 
 output OKA; 
 output OKB; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output OMG; 
 output OMH; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AHP ;
reg  AIA ;
reg  AIB ;
reg  AIC ;
reg  AID ;
reg  AIE ;
reg  AIF ;
reg  AIG ;
reg  AIH ;
reg  AII ;
reg  AIJ ;
reg  AIK ;
reg  AIL ;
reg  AIM ;
reg  AIN ;
reg  AIO ;
reg  AIP ;
reg  AJA ;
reg  AJB ;
reg  AJC ;
reg  AJD ;
reg  AJE ;
reg  AJF ;
reg  AJG ;
reg  AJH ;
reg  AJI ;
reg  AJJ ;
reg  AJK ;
reg  AJL ;
reg  AJM ;
reg  AJN ;
reg  AJO ;
reg  AJP ;
reg  AKA ;
reg  AKB ;
reg  AKC ;
reg  AKD ;
reg  AKE ;
reg  AKF ;
reg  AKG ;
reg  AKH ;
reg  AKI ;
reg  AKJ ;
reg  AKK ;
reg  AKL ;
reg  AKM ;
reg  AKN ;
reg  AKO ;
reg  AKP ;
reg  ALA ;
reg  ALB ;
reg  ALC ;
reg  ALD ;
reg  ALE ;
reg  ALF ;
reg  ALG ;
reg  ALH ;
reg  ALI ;
reg  ALJ ;
reg  ALK ;
reg  ALL ;
reg  ALM ;
reg  ALN ;
reg  ALO ;
reg  ALP ;
reg  AMA ;
reg  AMB ;
reg  AMC ;
reg  AMD ;
reg  AME ;
reg  AMF ;
reg  AMG ;
reg  AMH ;
reg  AMI ;
reg  AMJ ;
reg  AMK ;
reg  AML ;
reg  AMM ;
reg  AMN ;
reg  AMO ;
reg  AMP ;
reg  ANA ;
reg  ANB ;
reg  ANC ;
reg  AND ;
reg  ANE ;
reg  ANF ;
reg  ANG ;
reg  ANH ;
reg  ANI ;
reg  ANJ ;
reg  ANK ;
reg  ANL ;
reg  ANM ;
reg  ANN ;
reg  ANO ;
reg  ANP ;
reg  AOA ;
reg  AOB ;
reg  AOC ;
reg  AOD ;
reg  AOE ;
reg  AOF ;
reg  AOG ;
reg  AOH ;
reg  AOI ;
reg  AOJ ;
reg  AOK ;
reg  AOL ;
reg  AOM ;
reg  AON ;
reg  AOO ;
reg  AOP ;
reg  APA ;
reg  APB ;
reg  APC ;
reg  APD ;
reg  APE ;
reg  APF ;
reg  APG ;
reg  APH ;
reg  API ;
reg  APJ ;
reg  APK ;
reg  APL ;
reg  APM ;
reg  APN ;
reg  APO ;
reg  APP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CDA ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CGA ;
reg  CGB ;
reg  CGC ;
reg  CGD ;
reg  CHA ;
reg  CHB ;
reg  CHC ;
reg  CHD ;
reg  CIA ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DDA ;
reg  DDB ;
reg  DDC ;
reg  DDD ;
reg  DEA ;
reg  DEB ;
reg  DEC ;
reg  DED ;
reg  DFA ;
reg  DFB ;
reg  DFC ;
reg  DFD ;
reg  DGA ;
reg  DGB ;
reg  DGC ;
reg  DGD ;
reg  DHA ;
reg  DHB ;
reg  DHC ;
reg  DHD ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBH ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  ECD ;
reg  ECE ;
reg  ECF ;
reg  ECG ;
reg  ECH ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EEA ;
reg  EEB ;
reg  EEC ;
reg  EED ;
reg  EEE ;
reg  EEF ;
reg  EEG ;
reg  EEH ;
reg  EFA ;
reg  EFB ;
reg  EFC ;
reg  EFD ;
reg  EFE ;
reg  EFF ;
reg  EFG ;
reg  EFH ;
reg  EGA ;
reg  EGB ;
reg  EGC ;
reg  EGD ;
reg  EGE ;
reg  EGF ;
reg  EGG ;
reg  EGH ;
reg  EHA ;
reg  EHB ;
reg  EHC ;
reg  EHD ;
reg  EHE ;
reg  EHF ;
reg  EHG ;
reg  EHH ;
reg  eia ;
reg  eib ;
reg  eic ;
reg  eid ;
reg  eie ;
reg  eif ;
reg  eig ;
reg  eih ;
reg  eja ;
reg  ejb ;
reg  ejc ;
reg  ejd ;
reg  eje ;
reg  ejf ;
reg  ejg ;
reg  ejh ;
reg  eka ;
reg  ekb ;
reg  ekc ;
reg  ekd ;
reg  eke ;
reg  ekf ;
reg  ekg ;
reg  ekh ;
reg  ela ;
reg  elb ;
reg  elc ;
reg  eld ;
reg  ele ;
reg  elf ;
reg  elg ;
reg  elh ;
reg  ema ;
reg  emb ;
reg  emc ;
reg  emd ;
reg  eme ;
reg  emf ;
reg  emg ;
reg  emh ;
reg  ena ;
reg  enb ;
reg  enc ;
reg  end ;
reg  ene ;
reg  enf ;
reg  eng ;
reg  enh ;
reg  eoa ;
reg  eob ;
reg  eoc ;
reg  eod ;
reg  eoe ;
reg  eof ;
reg  eog ;
reg  eoh ;
reg  epa ;
reg  epb ;
reg  epc ;
reg  epd ;
reg  epe ;
reg  epf ;
reg  epg ;
reg  eph ;
reg  kaa ;
reg  kab ;
reg  kac ;
reg  kad ;
reg  kae ;
reg  kaf ;
reg  kag ;
reg  kah ;
reg  kba ;
reg  kbb ;
reg  kbc ;
reg  kbd ;
reg  kbe ;
reg  kbf ;
reg  kbg ;
reg  kbh ;
reg  kca ;
reg  kcb ;
reg  kcc ;
reg  kcd ;
reg  kce ;
reg  kcf ;
reg  kcg ;
reg  kch ;
reg  kda ;
reg  kdb ;
reg  kdc ;
reg  kdd ;
reg  kde ;
reg  kdf ;
reg  kdg ;
reg  kdh ;
reg  kea ;
reg  keb ;
reg  kec ;
reg  ked ;
reg  kee ;
reg  kef ;
reg  keg ;
reg  keh ;
reg  kfa ;
reg  kfb ;
reg  kfc ;
reg  kfd ;
reg  kfe ;
reg  kff ;
reg  kfg ;
reg  kfh ;
reg  kga ;
reg  kgb ;
reg  kgc ;
reg  kgd ;
reg  kge ;
reg  kgf ;
reg  kgg ;
reg  kgh ;
reg  kha ;
reg  khb ;
reg  khc ;
reg  khd ;
reg  khe ;
reg  khf ;
reg  khg ;
reg  khh ;
reg  laa ;
reg  lab ;
reg  lac ;
reg  lad ;
reg  lae ;
reg  laf ;
reg  maa ;
reg  mab ;
reg  mac ;
reg  mae ;
reg  maf ;
reg  mag ;
reg  naa ;
reg  nab ;
reg  nac ;
reg  nae ;
reg  naf ;
reg  nag ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  OHL ;
reg  OHM ;
reg  OHN ;
reg  OHO ;
reg  OHP ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OIJ ;
reg  oja ;
reg  ojb ;
reg  ojc ;
reg  ojd ;
reg  oje ;
reg  ojf ;
reg  OKA ;
reg  OKB ;
reg  ola ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  OME ;
reg  OMF ;
reg  OMG ;
reg  OMH ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  qca ;
reg  qcb ;
reg  qcc ;
reg  qcd ;
reg  qce ;
reg  qcf ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  qfe ;
reg  qff ;
reg  qfg ;
reg  QFH ;
reg  QKA ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  RAI ;
reg  RAJ ;
reg  RAK ;
reg  RAL ;
reg  RAM ;
reg  RAN ;
reg  RAO ;
reg  RAP ;
reg  RBA ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  RBH ;
reg  RBI ;
reg  RBJ ;
reg  RBK ;
reg  RBL ;
reg  RBM ;
reg  RBN ;
reg  RBO ;
reg  RBP ;
reg  RCA ;
reg  RCB ;
reg  RCC ;
reg  RCD ;
reg  RCE ;
reg  RCF ;
reg  RCG ;
reg  RCH ;
reg  RCI ;
reg  RCJ ;
reg  RCK ;
reg  RCL ;
reg  RCM ;
reg  RCN ;
reg  RCO ;
reg  RCP ;
reg  RDA ;
reg  RDB ;
reg  RDC ;
reg  RDD ;
reg  RDE ;
reg  RDF ;
reg  RDG ;
reg  RDH ;
reg  RDI ;
reg  RDJ ;
reg  RDK ;
reg  RDL ;
reg  RDM ;
reg  RDN ;
reg  RDO ;
reg  RDP ;
reg  RGA ;
reg  RGB ;
reg  RGC ;
reg  RGD ;
reg  RGE ;
reg  RGF ;
reg  RGG ;
reg  RGH ;
reg  RGI ;
reg  RGJ ;
reg  RGK ;
reg  RGL ;
reg  RGM ;
reg  RGN ;
reg  RGO ;
reg  RGP ;
reg  RHA ;
reg  RHB ;
reg  RHC ;
reg  RHD ;
reg  RHE ;
reg  RHF ;
reg  RHG ;
reg  RHH ;
reg  RHI ;
reg  RHJ ;
reg  RHK ;
reg  RHL ;
reg  RHM ;
reg  RHN ;
reg  RHO ;
reg  RHP ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  SAD ;
reg  SAE ;
reg  SAF ;
reg  SAG ;
reg  SAH ;
reg  SAI ;
reg  SAJ ;
reg  SAK ;
reg  SAL ;
reg  SAM ;
reg  SAN ;
reg  SAO ;
reg  SAP ;
reg  SBA ;
reg  SBB ;
reg  SBC ;
reg  SBD ;
reg  SBE ;
reg  SBF ;
reg  SBG ;
reg  SBH ;
reg  SBI ;
reg  SBJ ;
reg  SBK ;
reg  SBL ;
reg  SBM ;
reg  SBN ;
reg  SBO ;
reg  SBP ;
reg  SCM ;
reg  SCN ;
reg  SCO ;
reg  SCP ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TAI ;
reg  TAJ ;
reg  TAK ;
reg  TAL ;
reg  TAM ;
reg  TAN ;
reg  TAO ;
reg  TAP ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TIA ;
reg  TIB ;
reg  TIC ;
reg  TID ;
reg  TIE ;
reg  TIF ;
reg  TIG ;
reg  TIH ;
reg  TJA ;
reg  TJB ;
reg  TJC ;
reg  TJD ;
reg  TJE ;
reg  TJF ;
reg  TJG ;
reg  TJH ;
reg  TKA ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  TKE ;
reg  TKF ;
reg  TKG ;
reg  TKH ;
reg  TKI ;
reg  TKJ ;
reg  TKK ;
reg  TKL ;
reg  TKM ;
reg  TKN ;
reg  TKO ;
reg  TKP ;
reg  TLA ;
reg  TLB ;
reg  TLC ;
reg  TLD ;
reg  TLE ;
reg  TLF ;
reg  TLG ;
reg  TLH ;
reg  TLI ;
reg  TLJ ;
reg  TLK ;
reg  TLL ;
reg  TLM ;
reg  TLN ;
reg  TLO ;
reg  TLP ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TMD ;
reg  TME ;
reg  TMF ;
reg  TMG ;
reg  TMH ;
reg  TMI ;
reg  TMJ ;
reg  TMK ;
reg  TML ;
reg  TMM ;
reg  TMN ;
reg  TMO ;
reg  TMP ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  ahp ;
wire  aia ;
wire  aib ;
wire  aic ;
wire  aid ;
wire  aie ;
wire  aif ;
wire  aig ;
wire  aih ;
wire  aii ;
wire  aij ;
wire  aik ;
wire  ail ;
wire  aim ;
wire  ain ;
wire  aio ;
wire  aip ;
wire  aja ;
wire  ajb ;
wire  ajc ;
wire  ajd ;
wire  aje ;
wire  ajf ;
wire  ajg ;
wire  ajh ;
wire  aji ;
wire  ajj ;
wire  ajk ;
wire  ajl ;
wire  ajm ;
wire  ajn ;
wire  ajo ;
wire  ajp ;
wire  aka ;
wire  akb ;
wire  akc ;
wire  akd ;
wire  ake ;
wire  akf ;
wire  akg ;
wire  akh ;
wire  aki ;
wire  akj ;
wire  akk ;
wire  akl ;
wire  akm ;
wire  akn ;
wire  ako ;
wire  akp ;
wire  ala ;
wire  alb ;
wire  alc ;
wire  ald ;
wire  ale ;
wire  alf ;
wire  alg ;
wire  alh ;
wire  ali ;
wire  alj ;
wire  alk ;
wire  all ;
wire  alm ;
wire  aln ;
wire  alo ;
wire  alp ;
wire  ama ;
wire  amb ;
wire  amc ;
wire  amd ;
wire  ame ;
wire  amf ;
wire  amg ;
wire  amh ;
wire  ami ;
wire  amj ;
wire  amk ;
wire  aml ;
wire  amm ;
wire  amn ;
wire  amo ;
wire  amp ;
wire  ana ;
wire  anb ;
wire  anc ;
wire  and ;
wire  ane ;
wire  anf ;
wire  ang ;
wire  anh ;
wire  ani ;
wire  anj ;
wire  ank ;
wire  anl ;
wire  anm ;
wire  ann ;
wire  ano ;
wire  anp ;
wire  aoa ;
wire  aob ;
wire  aoc ;
wire  aod ;
wire  aoe ;
wire  aof ;
wire  aog ;
wire  aoh ;
wire  aoi ;
wire  aoj ;
wire  aok ;
wire  aol ;
wire  aom ;
wire  aon ;
wire  aoo ;
wire  aop ;
wire  apa ;
wire  apb ;
wire  apc ;
wire  apd ;
wire  ape ;
wire  apf ;
wire  apg ;
wire  aph ;
wire  api ;
wire  apj ;
wire  apk ;
wire  apl ;
wire  apm ;
wire  apn ;
wire  apo ;
wire  app ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cda ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cga ;
wire  cgb ;
wire  cgc ;
wire  cgd ;
wire  cha ;
wire  chb ;
wire  chc ;
wire  chd ;
wire  cia ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dda ;
wire  ddb ;
wire  ddc ;
wire  ddd ;
wire  dea ;
wire  deb ;
wire  dec ;
wire  ded ;
wire  dfa ;
wire  dfb ;
wire  dfc ;
wire  dfd ;
wire  dga ;
wire  dgb ;
wire  dgc ;
wire  dgd ;
wire  dha ;
wire  dhb ;
wire  dhc ;
wire  dhd ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebh ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  ecd ;
wire  ece ;
wire  ecf ;
wire  ecg ;
wire  ech ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  eea ;
wire  eeb ;
wire  eec ;
wire  eed ;
wire  eee ;
wire  eef ;
wire  eeg ;
wire  eeh ;
wire  efa ;
wire  efb ;
wire  efc ;
wire  efd ;
wire  efe ;
wire  eff ;
wire  efg ;
wire  efh ;
wire  ega ;
wire  egb ;
wire  egc ;
wire  egd ;
wire  ege ;
wire  egf ;
wire  egg ;
wire  egh ;
wire  eha ;
wire  ehb ;
wire  ehc ;
wire  ehd ;
wire  ehe ;
wire  ehf ;
wire  ehg ;
wire  ehh ;
wire  EIA ;
wire  EIB ;
wire  EIC ;
wire  EID ;
wire  EIE ;
wire  EIF ;
wire  EIG ;
wire  EIH ;
wire  EJA ;
wire  EJB ;
wire  EJC ;
wire  EJD ;
wire  EJE ;
wire  EJF ;
wire  EJG ;
wire  EJH ;
wire  EKA ;
wire  EKB ;
wire  EKC ;
wire  EKD ;
wire  EKE ;
wire  EKF ;
wire  EKG ;
wire  EKH ;
wire  ELA ;
wire  ELB ;
wire  ELC ;
wire  ELD ;
wire  ELE ;
wire  ELF ;
wire  ELG ;
wire  ELH ;
wire  EMA ;
wire  EMB ;
wire  EMC ;
wire  EMD ;
wire  EME ;
wire  EMF ;
wire  EMG ;
wire  EMH ;
wire  ENA ;
wire  ENB ;
wire  ENC ;
wire  END ;
wire  ENE ;
wire  ENF ;
wire  ENG ;
wire  ENH ;
wire  EOA ;
wire  EOB ;
wire  EOC ;
wire  EOD ;
wire  EOE ;
wire  EOF ;
wire  EOG ;
wire  EOH ;
wire  EPA ;
wire  EPB ;
wire  EPC ;
wire  EPD ;
wire  EPE ;
wire  EPF ;
wire  EPG ;
wire  EPH ;
wire  FAA ;
wire  FAB ;
wire  FAC ;
wire  FAD ;
wire  FAE ;
wire  FAF ;
wire  FAG ;
wire  FAH ;
wire  FAI ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gbf ;
wire  GBF ;
wire  gbg ;
wire  GBG ;
wire  gbh ;
wire  GBH ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  haa ;
wire  HAA ;
wire  hab ;
wire  HAB ;
wire  hac ;
wire  HAC ;
wire  had ;
wire  HAD ;
wire  hae ;
wire  HAE ;
wire  hba ;
wire  HBA ;
wire  hbb ;
wire  HBB ;
wire  hbc ;
wire  HBC ;
wire  hbd ;
wire  HBD ;
wire  hbe ;
wire  HBE ;
wire  hca ;
wire  HCA ;
wire  hcb ;
wire  HCB ;
wire  hcc ;
wire  HCC ;
wire  hcd ;
wire  HCD ;
wire  hce ;
wire  HCE ;
wire  hda ;
wire  HDA ;
wire  hdb ;
wire  HDB ;
wire  hdc ;
wire  HDC ;
wire  hdd ;
wire  HDD ;
wire  hde ;
wire  HDE ;
wire  hea ;
wire  HEA ;
wire  heb ;
wire  HEB ;
wire  hec ;
wire  HEC ;
wire  hed ;
wire  HED ;
wire  hee ;
wire  HEE ;
wire  hfa ;
wire  HFA ;
wire  hfb ;
wire  HFB ;
wire  hfc ;
wire  HFC ;
wire  hfd ;
wire  HFD ;
wire  hfe ;
wire  HFE ;
wire  hga ;
wire  HGA ;
wire  hgb ;
wire  HGB ;
wire  hgc ;
wire  HGC ;
wire  hgd ;
wire  HGD ;
wire  hge ;
wire  HGE ;
wire  hha ;
wire  HHA ;
wire  hhb ;
wire  HHB ;
wire  hhc ;
wire  HHC ;
wire  hhd ;
wire  HHD ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iff ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  ihm ;
wire  ihn ;
wire  iho ;
wire  ihp ;
wire  iia ;
wire  iib ;
wire  iic ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  ika ;
wire  ikb ;
wire  ila ;
wire  ima ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jbo ;
wire  JBO ;
wire  jbp ;
wire  JBP ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jci ;
wire  JCI ;
wire  jcj ;
wire  JCJ ;
wire  jck ;
wire  JCK ;
wire  jcl ;
wire  JCL ;
wire  jcm ;
wire  JCM ;
wire  jcn ;
wire  JCN ;
wire  jco ;
wire  JCO ;
wire  jcp ;
wire  JCP ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jdp ;
wire  JDP ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jei ;
wire  JEI ;
wire  jej ;
wire  JEJ ;
wire  jek ;
wire  JEK ;
wire  jel ;
wire  JEL ;
wire  jem ;
wire  JEM ;
wire  jen ;
wire  JEN ;
wire  jeo ;
wire  JEO ;
wire  jep ;
wire  JEP ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jfi ;
wire  JFI ;
wire  jfj ;
wire  JFJ ;
wire  jfk ;
wire  JFK ;
wire  jfl ;
wire  JFL ;
wire  jfm ;
wire  JFM ;
wire  jfn ;
wire  JFN ;
wire  jfo ;
wire  JFO ;
wire  jfp ;
wire  JFP ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgh ;
wire  JGH ;
wire  jgi ;
wire  JGI ;
wire  jgj ;
wire  JGJ ;
wire  jgk ;
wire  JGK ;
wire  jgl ;
wire  JGL ;
wire  jgm ;
wire  JGM ;
wire  jgn ;
wire  JGN ;
wire  jgo ;
wire  JGO ;
wire  jgp ;
wire  JGP ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jhi ;
wire  JHI ;
wire  jhj ;
wire  JHJ ;
wire  jhk ;
wire  JHK ;
wire  jhl ;
wire  JHL ;
wire  jhm ;
wire  JHM ;
wire  jhn ;
wire  JHN ;
wire  jho ;
wire  JHO ;
wire  jhp ;
wire  JHP ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jie ;
wire  JIE ;
wire  jif ;
wire  JIF ;
wire  jig ;
wire  JIG ;
wire  jih ;
wire  JIH ;
wire  KAA ;
wire  KAB ;
wire  KAC ;
wire  KAD ;
wire  KAE ;
wire  KAF ;
wire  KAG ;
wire  KAH ;
wire  KBA ;
wire  KBB ;
wire  KBC ;
wire  KBD ;
wire  KBE ;
wire  KBF ;
wire  KBG ;
wire  KBH ;
wire  KCA ;
wire  KCB ;
wire  KCC ;
wire  KCD ;
wire  KCE ;
wire  KCF ;
wire  KCG ;
wire  KCH ;
wire  KDA ;
wire  KDB ;
wire  KDC ;
wire  KDD ;
wire  KDE ;
wire  KDF ;
wire  KDG ;
wire  KDH ;
wire  KEA ;
wire  KEB ;
wire  KEC ;
wire  KED ;
wire  KEE ;
wire  KEF ;
wire  KEG ;
wire  KEH ;
wire  KFA ;
wire  KFB ;
wire  KFC ;
wire  KFD ;
wire  KFE ;
wire  KFF ;
wire  KFG ;
wire  KFH ;
wire  KGA ;
wire  KGB ;
wire  KGC ;
wire  KGD ;
wire  KGE ;
wire  KGF ;
wire  KGG ;
wire  KGH ;
wire  KHA ;
wire  KHB ;
wire  KHC ;
wire  KHD ;
wire  KHE ;
wire  KHF ;
wire  KHG ;
wire  KHH ;
wire  LAA ;
wire  LAB ;
wire  LAC ;
wire  LAD ;
wire  LAE ;
wire  LAF ;
wire  MAA ;
wire  MAB ;
wire  MAC ;
wire  MAE ;
wire  MAF ;
wire  MAG ;
wire  NAA ;
wire  NAB ;
wire  NAC ;
wire  NAE ;
wire  NAF ;
wire  NAG ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  ohl ;
wire  ohm ;
wire  ohn ;
wire  oho ;
wire  ohp ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oij ;
wire  OJA ;
wire  OJB ;
wire  OJC ;
wire  OJD ;
wire  OJE ;
wire  OJF ;
wire  oka ;
wire  okb ;
wire  OLA ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  ome ;
wire  omf ;
wire  omg ;
wire  omh ;
wire  paa ;
wire  PAA ;
wire  pab ;
wire  PAB ;
wire  pac ;
wire  PAC ;
wire  pad ;
wire  PAD ;
wire  pae ;
wire  PAE ;
wire  paf ;
wire  PAF ;
wire  pag ;
wire  PAG ;
wire  pah ;
wire  PAH ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  QCA ;
wire  QCB ;
wire  QCC ;
wire  QCD ;
wire  QCE ;
wire  QCF ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  QFE ;
wire  QFF ;
wire  QFG ;
wire  qfh ;
wire  qha ;
wire  QHA ;
wire  qhb ;
wire  QHB ;
wire  qhc ;
wire  QHC ;
wire  qhd ;
wire  QHD ;
wire  qhe ;
wire  QHE ;
wire  qhf ;
wire  QHF ;
wire  qhg ;
wire  QHG ;
wire  qhh ;
wire  QHH ;
wire  qia ;
wire  QIA ;
wire  qib ;
wire  QIB ;
wire  qic ;
wire  QIC ;
wire  qid ;
wire  QID ;
wire  qie ;
wire  QIE ;
wire  qif ;
wire  QIF ;
wire  qig ;
wire  QIG ;
wire  qih ;
wire  QIH ;
wire  qja ;
wire  QJA ;
wire  qjb ;
wire  QJB ;
wire  qjc ;
wire  QJC ;
wire  qjd ;
wire  QJD ;
wire  qje ;
wire  QJE ;
wire  qjf ;
wire  QJF ;
wire  qjg ;
wire  QJG ;
wire  qjh ;
wire  QJH ;
wire  qji ;
wire  QJI ;
wire  qjj ;
wire  QJJ ;
wire  qjk ;
wire  QJK ;
wire  qjl ;
wire  QJL ;
wire  qka ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  rai ;
wire  raj ;
wire  rak ;
wire  ral ;
wire  ram ;
wire  ran ;
wire  rao ;
wire  rap ;
wire  rba ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  rbh ;
wire  rbi ;
wire  rbj ;
wire  rbk ;
wire  rbl ;
wire  rbm ;
wire  rbn ;
wire  rbo ;
wire  rbp ;
wire  rca ;
wire  rcb ;
wire  rcc ;
wire  rcd ;
wire  rce ;
wire  rcf ;
wire  rcg ;
wire  rch ;
wire  rci ;
wire  rcj ;
wire  rck ;
wire  rcl ;
wire  rcm ;
wire  rcn ;
wire  rco ;
wire  rcp ;
wire  rda ;
wire  rdb ;
wire  rdc ;
wire  rdd ;
wire  rde ;
wire  rdf ;
wire  rdg ;
wire  rdh ;
wire  rdi ;
wire  rdj ;
wire  rdk ;
wire  rdl ;
wire  rdm ;
wire  rdn ;
wire  rdo ;
wire  rdp ;
wire  rea ;
wire  REA ;
wire  reb ;
wire  REB ;
wire  rec ;
wire  REC ;
wire  red ;
wire  RED ;
wire  ree ;
wire  REE ;
wire  ref ;
wire  REF ;
wire  reg ;
wire  REG ;
wire  reh ;
wire  REH ;
wire  rei ;
wire  REI ;
wire  rej ;
wire  REJ ;
wire  rek ;
wire  REK ;
wire  rel ;
wire  REL ;
wire  rem ;
wire  REM ;
wire  ren ;
wire  REN ;
wire  reo ;
wire  REO ;
wire  rep ;
wire  REP ;
wire  rfa ;
wire  RFA ;
wire  rfb ;
wire  RFB ;
wire  rfc ;
wire  RFC ;
wire  rfd ;
wire  RFD ;
wire  rfe ;
wire  RFE ;
wire  rff ;
wire  RFF ;
wire  rfg ;
wire  RFG ;
wire  rfh ;
wire  RFH ;
wire  rfi ;
wire  RFI ;
wire  rfj ;
wire  RFJ ;
wire  rfk ;
wire  RFK ;
wire  rfl ;
wire  RFL ;
wire  rfm ;
wire  RFM ;
wire  rfn ;
wire  RFN ;
wire  rfo ;
wire  RFO ;
wire  rfp ;
wire  RFP ;
wire  rga ;
wire  rgb ;
wire  rgc ;
wire  rgd ;
wire  rge ;
wire  rgf ;
wire  rgg ;
wire  rgh ;
wire  rgi ;
wire  rgj ;
wire  rgk ;
wire  rgl ;
wire  rgm ;
wire  rgn ;
wire  rgo ;
wire  rgp ;
wire  rha ;
wire  rhb ;
wire  rhc ;
wire  rhd ;
wire  rhe ;
wire  rhf ;
wire  rhg ;
wire  rhh ;
wire  rhi ;
wire  rhj ;
wire  rhk ;
wire  rhl ;
wire  rhm ;
wire  rhn ;
wire  rho ;
wire  rhp ;
wire  ria ;
wire  RIA ;
wire  rib ;
wire  RIB ;
wire  ric ;
wire  RIC ;
wire  rid ;
wire  RID ;
wire  rie ;
wire  RIE ;
wire  rif ;
wire  RIF ;
wire  rig ;
wire  RIG ;
wire  rih ;
wire  RIH ;
wire  rii ;
wire  RII ;
wire  rij ;
wire  RIJ ;
wire  rik ;
wire  RIK ;
wire  ril ;
wire  RIL ;
wire  rim ;
wire  RIM ;
wire  rin ;
wire  RIN ;
wire  rio ;
wire  RIO ;
wire  rip ;
wire  RIP ;
wire  rja ;
wire  RJA ;
wire  rjb ;
wire  RJB ;
wire  rjc ;
wire  RJC ;
wire  rjd ;
wire  RJD ;
wire  rje ;
wire  RJE ;
wire  rjf ;
wire  RJF ;
wire  rjg ;
wire  RJG ;
wire  rjh ;
wire  RJH ;
wire  rji ;
wire  RJI ;
wire  rjj ;
wire  RJJ ;
wire  rjk ;
wire  RJK ;
wire  rjl ;
wire  RJL ;
wire  rjm ;
wire  RJM ;
wire  rjn ;
wire  RJN ;
wire  rjo ;
wire  RJO ;
wire  rjp ;
wire  RJP ;
wire  saa ;
wire  sab ;
wire  sac ;
wire  sad ;
wire  sae ;
wire  saf ;
wire  sag ;
wire  sah ;
wire  sai ;
wire  saj ;
wire  sak ;
wire  sal ;
wire  sam ;
wire  san ;
wire  sao ;
wire  sap ;
wire  sba ;
wire  sbb ;
wire  sbc ;
wire  sbd ;
wire  sbe ;
wire  sbf ;
wire  sbg ;
wire  sbh ;
wire  sbi ;
wire  sbj ;
wire  sbk ;
wire  sbl ;
wire  sbm ;
wire  sbn ;
wire  sbo ;
wire  sbp ;
wire  scm ;
wire  scn ;
wire  sco ;
wire  scp ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tai ;
wire  taj ;
wire  tak ;
wire  tal ;
wire  tam ;
wire  tan ;
wire  tao ;
wire  tap ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tcg ;
wire  TCG ;
wire  tch ;
wire  TCH ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tde ;
wire  TDE ;
wire  tdf ;
wire  TDF ;
wire  tdg ;
wire  TDG ;
wire  tdh ;
wire  TDH ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  teg ;
wire  TEG ;
wire  teh ;
wire  TEH ;
wire  tfa ;
wire  TFA ;
wire  tfb ;
wire  TFB ;
wire  tfc ;
wire  TFC ;
wire  tfd ;
wire  TFD ;
wire  tfe ;
wire  TFE ;
wire  tff ;
wire  TFF ;
wire  tfg ;
wire  TFG ;
wire  tfh ;
wire  TFH ;
wire  tia ;
wire  tib ;
wire  tic ;
wire  tid ;
wire  tie ;
wire  tif ;
wire  tig ;
wire  tih ;
wire  tja ;
wire  tjb ;
wire  tjc ;
wire  tjd ;
wire  tje ;
wire  tjf ;
wire  tjg ;
wire  tjh ;
wire  tka ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  tke ;
wire  tkf ;
wire  tkg ;
wire  tkh ;
wire  tki ;
wire  tkj ;
wire  tkk ;
wire  tkl ;
wire  tkm ;
wire  tkn ;
wire  tko ;
wire  tkp ;
wire  tla ;
wire  tlb ;
wire  tlc ;
wire  tld ;
wire  tle ;
wire  tlf ;
wire  tlg ;
wire  tlh ;
wire  tli ;
wire  tlj ;
wire  tlk ;
wire  tll ;
wire  tlm ;
wire  tln ;
wire  tlo ;
wire  tlp ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tmd ;
wire  tme ;
wire  tmf ;
wire  tmg ;
wire  tmh ;
wire  tmi ;
wire  tmj ;
wire  tmk ;
wire  tml ;
wire  tmm ;
wire  tmn ;
wire  tmo ;
wire  tmp ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign GAB =  CAA  ; 
assign gab = ~GAB;  //complement 
assign GAC =  CAA & DAB  |  CAB  ; 
assign gac = ~GAC;  //complement 
assign caa = ~CAA;  //complement 
assign daa = ~DAA;  //complement 
assign GAD =  CAA & DAB & DAC  |  CAB & DAC  |  CAC  ; 
assign gad = ~GAD;  //complement 
assign cab = ~CAB;  //complement 
assign dab = ~DAB;  //complement 
assign KAA = ~kaa;  //complement 
assign KAE = ~kae;  //complement 
assign GAE =  CAA & DAB & DAC & DAD  |  CAB & DAC & DAD  |  CAC & DAD  |  CAD  ; 
assign gae = ~GAE;  //complement 
assign KAB = ~kab;  //complement 
assign KAF = ~kaf;  //complement 
assign MAA = ~maa;  //complement 
assign NAA = ~naa;  //complement 
assign KEB = ~keb;  //complement 
assign KEF = ~kef;  //complement 
assign MAE = ~mae;  //complement 
assign NAE = ~nae;  //complement 
assign KEA = ~kea;  //complement 
assign KEE = ~kee;  //complement 
assign GEE =  CEA & DEB & DEC & DED  |  CEB & DEC & DED  |  CEC & DED  |  CED  ; 
assign gee = ~GEE;  //complement 
assign GED =  CEA & DEB & DEC  |  CEB & DEC  |  CEC  ; 
assign ged = ~GED;  //complement 
assign cea = ~CEA;  //complement 
assign dea = ~DEA;  //complement 
assign GEB =  CEA  ; 
assign geb = ~GEB;  //complement 
assign GEC =  CEA & DEB  |  CEB  ; 
assign gec = ~GEC;  //complement 
assign ceb = ~CEB;  //complement 
assign deb = ~DEB;  //complement 
assign baa = ~BAA;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign JAA =  AAA & EAA  |  ABA & EBA  |  ACA & ECA  |  ADA & EDA  |  CIA  ;
assign jaa = ~JAA;  //complement 
assign bab = ~BAB;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign eaa = ~EAA;  //complement 
assign eba = ~EBA;  //complement 
assign eca = ~ECA;  //complement 
assign eda = ~EDA;  //complement 
assign raa = ~RAA;  //complement 
assign rab = ~RAB;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign QJA = QFE; 
assign qja = ~QJA; //complement 
assign QJB = QFE; 
assign qjb = ~QJB;  //complement 
assign qjc = qfe; 
assign QJC = ~qjc;  //complement 
assign qjd = qfe; 
assign QJD = ~qjd;  //complement 
assign REA = RAA; 
assign rea = ~REA; //complement 
assign REB = RAB; 
assign reb = ~REB;  //complement 
assign RIA = RAA; 
assign ria = ~RIA;  //complement 
assign RIB = RAB; 
assign rib = ~RIB;  //complement 
assign tad = ~TAD;  //complement 
assign tal = ~TAL;  //complement 
assign tkd = ~TKD;  //complement 
assign tkl = ~TKL;  //complement 
assign aga = ~AGA;  //complement 
assign agb = ~AGB;  //complement 
assign eea = ~EEA;  //complement 
assign efa = ~EFA;  //complement 
assign ega = ~EGA;  //complement 
assign eha = ~EHA;  //complement 
assign RFA = RBA; 
assign rfa = ~RFA; //complement 
assign RFB = RBB; 
assign rfb = ~RFB;  //complement 
assign RJA = RBA; 
assign rja = ~RJA;  //complement 
assign RJB = RBB; 
assign rjb = ~RJB;  //complement 
assign tah = ~TAH;  //complement 
assign tap = ~TAP;  //complement 
assign tkh = ~TKH;  //complement 
assign tkp = ~TKP;  //complement 
assign aia = ~AIA;  //complement 
assign aib = ~AIB;  //complement 
assign EIA = ~eia;  //complement 
assign EJA = ~eja;  //complement 
assign EKA = ~eka;  //complement 
assign rba = ~RBA;  //complement 
assign rbb = ~RBB;  //complement 
assign aka = ~AKA;  //complement 
assign akb = ~AKB;  //complement 
assign ELA = ~ela;  //complement 
assign EPA = ~epa;  //complement 
assign bea = ~BEA;  //complement 
assign ama = ~AMA;  //complement 
assign amb = ~AMB;  //complement 
assign EMA = ~ema;  //complement 
assign ENA = ~ena;  //complement 
assign EOA = ~eoa;  //complement 
assign beb = ~BEB;  //complement 
assign aoa = ~AOA;  //complement 
assign aob = ~AOB;  //complement 
assign JEA =  AAA & EAA  |  ABA & EBA  |  ACA & ECA  |  ADA & EDA  ; 
assign jea = ~JEA;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign rca = ~RCA;  //complement 
assign rga = ~RGA;  //complement 
assign LAA = ~laa;  //complement 
assign OJA = ~oja;  //complement 
assign JAB =  AAB & EAA  |  ABB & EBA  |  ACB & ECA  |  ADB & EDA  ; 
assign jab = ~JAB;  //complement 
assign JEB =  AAB & EAA  |  ABB & EBA  |  ACB & ECA  |  ADB & EDA  ; 
assign jeb = ~JEB; //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign rcb = ~RCB;  //complement 
assign rgb = ~RGB;  //complement 
assign LAB = ~lab;  //complement 
assign OJB = ~ojb;  //complement 
assign JBA =  AEA & EEA  |  AFA & EFA  |  AGA & EGA  |  AHA & EHA  ; 
assign jba = ~JBA;  //complement 
assign JFA =  AEA & EEA  |  AFA & EFA  |  AGA & EGA  |  AHA & EHA  ; 
assign jfa = ~JFA; //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign oga = ~OGA;  //complement 
assign oia = ~OIA;  //complement 
assign saa = ~SAA;  //complement 
assign oaa = ~OAA;  //complement 
assign oca = ~OCA;  //complement 
assign oea = ~OEA;  //complement 
assign JBB =  AEB & EEA  |  AFB & EFA  |  AGB & EGA  |  AHB & EHA  ; 
assign jbb = ~JBB;  //complement 
assign JFB =  AEB & EEA  |  AFB & EFA  |  AGB & EGA  |  AHB & EHA  ; 
assign jfb = ~JFB; //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign ogb = ~OGB;  //complement 
assign oib = ~OIB;  //complement 
assign sab = ~SAB;  //complement 
assign oab = ~OAB;  //complement 
assign ocb = ~OCB;  //complement 
assign oeb = ~OEB;  //complement 
assign JCA =  AIA & EIA  |  AJA & EJA  |  AKA & EKA  |  ALA & ELA  ; 
assign jca = ~JCA;  //complement 
assign JGA =  AIA & EIA  |  AJA & EJA  |  AKA & EKA  |  ALA & ELA  ; 
assign jga = ~JGA; //complement 
assign aja = ~AJA;  //complement 
assign ajb = ~AJB;  //complement 
assign oha = ~OHA;  //complement 
assign sba = ~SBA;  //complement 
assign oba = ~OBA;  //complement 
assign oda = ~ODA;  //complement 
assign ofa = ~OFA;  //complement 
assign JCB =  AIB & EIA  |  AJB & EJA  |  AKB & EKA  |  ALB & ELA  ; 
assign jcb = ~JCB;  //complement 
assign JGB =  AIB & EIA  |  AJB & EJA  |  AKB & EKA  |  ALB & ELA  ; 
assign jgb = ~JGB; //complement 
assign ala = ~ALA;  //complement 
assign alb = ~ALB;  //complement 
assign ohb = ~OHB;  //complement 
assign sbb = ~SBB;  //complement 
assign obb = ~OBB;  //complement 
assign odb = ~ODB;  //complement 
assign ofb = ~OFB;  //complement 
assign JDA =  AMA & EMA  |  ANA & ENA  |  AOA & EOA  |  APA & EPA  ; 
assign jda = ~JDA;  //complement 
assign JHA =  AMA & EMA  |  ANA & ENA  |  AOA & EOA  |  APA & EPA  ; 
assign jha = ~JHA; //complement 
assign ana = ~ANA;  //complement 
assign anb = ~ANB;  //complement 
assign rda = ~RDA;  //complement 
assign rha = ~RHA;  //complement 
assign cia = ~CIA;  //complement 
assign JDB =  AMB & EMA  |  ANB & ENA  |  AOB & EOA  |  APB & EPA  ; 
assign jdb = ~JDB;  //complement 
assign JHB =  AMB & EMA  |  ANB & ENA  |  AOB & EOA  |  APB & EPA  ; 
assign jhb = ~JHB; //complement 
assign apa = ~APA;  //complement 
assign apb = ~APB;  //complement 
assign rdb = ~RDB;  //complement 
assign rhb = ~RHB;  //complement 
assign gaf =  daa  ; 
assign GAF = ~gaf;  //complement 
assign gag =  daa & cab  |  dab  ; 
assign GAG = ~gag;  //complement 
assign cac = ~CAC;  //complement 
assign dac = ~DAC;  //complement 
assign gah =  daa & cab & cac  |  dab & cac  |  dac  ; 
assign GAH = ~gah;  //complement 
assign cad = ~CAD;  //complement 
assign dad = ~DAD;  //complement 
assign KAC = ~kac;  //complement 
assign KAG = ~kag;  //complement 
assign HAA =  DAA & caa  ; 
assign haa = ~HAA;  //complement 
assign HAB =  DAB & cab  ; 
assign hab = ~HAB;  //complement 
assign HAC =  DAC & cac  ; 
assign hac = ~HAC;  //complement 
assign PAA =  QAE  ; 
assign paa = ~PAA;  //complement 
assign KAD = ~kad;  //complement 
assign KAH = ~kah;  //complement 
assign HAD =  DAD & cad  ; 
assign had = ~HAD;  //complement  
assign HAE =  DAA & DAB & DAC & DAD  ; 
assign hae = ~HAE;  //complement 
assign KED = ~ked;  //complement 
assign KEH = ~keh;  //complement 
assign HED =  DED & ced  ; 
assign hed = ~HED;  //complement  
assign HEE =  DEA & DEB & DEC & DED  ; 
assign hee = ~HEE;  //complement 
assign tag = ~TAG;  //complement 
assign tao = ~TAO;  //complement 
assign tkg = ~TKG;  //complement 
assign tko = ~TKO;  //complement 
assign KEC = ~kec;  //complement 
assign KEG = ~keg;  //complement 
assign HEA =  DEA & cea  ; 
assign hea = ~HEA;  //complement 
assign HEB =  DEB & ceb  ; 
assign heb = ~HEB;  //complement 
assign HEC =  DEC & cec  ; 
assign hec = ~HEC;  //complement 
assign PAE =  QAF  ; 
assign pae = ~PAE;  //complement 
assign geh =  dea & ceb & cec  |  deb & cec  |  dec  ; 
assign GEH = ~geh;  //complement 
assign cec = ~CEC;  //complement 
assign dec = ~DEC;  //complement 
assign gef =  dea  ; 
assign GEF = ~gef;  //complement 
assign geg =  dea & ceb  |  deb  ; 
assign GEG = ~geg;  //complement 
assign ced = ~CED;  //complement 
assign ded = ~DED;  //complement 
assign bac = ~BAC;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign bad = ~BAD;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign eab = ~EAB;  //complement 
assign ebb = ~EBB;  //complement 
assign ecb = ~ECB;  //complement 
assign edb = ~EDB;  //complement 
assign rac = ~RAC;  //complement 
assign rad = ~RAD;  //complement 
assign aec = ~AEC;  //complement 
assign aed = ~AED;  //complement 
assign QJE = QFF; 
assign qje = ~QJE; //complement 
assign QJF = QFF; 
assign qjf = ~QJF;  //complement 
assign qjg = qff; 
assign QJG = ~qjg;  //complement 
assign qjh = qff; 
assign QJH = ~qjh;  //complement 
assign REC = RAC; 
assign rec = ~REC; //complement 
assign RED = RAD; 
assign red = ~RED;  //complement 
assign RIC = RAC; 
assign ric = ~RIC;  //complement 
assign RID = RAD; 
assign rid = ~RID;  //complement 
assign tac = ~TAC;  //complement 
assign tak = ~TAK;  //complement 
assign tkc = ~TKC;  //complement 
assign tkk = ~TKK;  //complement 
assign agc = ~AGC;  //complement 
assign agd = ~AGD;  //complement 
assign eeb = ~EEB;  //complement 
assign efb = ~EFB;  //complement 
assign egb = ~EGB;  //complement 
assign ehb = ~EHB;  //complement 
assign RFC = RBC; 
assign rfc = ~RFC; //complement 
assign RFD = RBD; 
assign rfd = ~RFD;  //complement 
assign RJC = RBC; 
assign rjc = ~RJC;  //complement 
assign RJD = RBD; 
assign rjd = ~RJD;  //complement 
assign QJI = QFG; 
assign qji = ~QJI; //complement 
assign QJJ = QFG; 
assign qjj = ~QJJ;  //complement 
assign qjk = qfg; 
assign QJK = ~qjk;  //complement 
assign qjl = qfg; 
assign QJL = ~qjl;  //complement 
assign aic = ~AIC;  //complement 
assign aid = ~AID;  //complement 
assign EIB = ~eib;  //complement 
assign EJB = ~ejb;  //complement 
assign EKB = ~ekb;  //complement 
assign rbc = ~RBC;  //complement 
assign rbd = ~RBD;  //complement 
assign akc = ~AKC;  //complement 
assign akd = ~AKD;  //complement 
assign ELB = ~elb;  //complement 
assign EPB = ~epb;  //complement 
assign bec = ~BEC;  //complement 
assign amc = ~AMC;  //complement 
assign amd = ~AMD;  //complement 
assign EMB = ~emb;  //complement 
assign ENB = ~enb;  //complement 
assign EOB = ~eob;  //complement 
assign bed = ~BED;  //complement 
assign aoc = ~AOC;  //complement 
assign aod = ~AOD;  //complement 
assign JAC =  AAC & EAB  |  ABC & EBB  |  ACC & ECB  |  ADC & EDB  ; 
assign jac = ~JAC;  //complement 
assign JEC =  AAC & EAB  |  ABC & EBB  |  ACC & ECB  |  ADC & EDB  ; 
assign jec = ~JEC; //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign rcc = ~RCC;  //complement 
assign rgc = ~RGC;  //complement 
assign LAC = ~lac;  //complement 
assign OJC = ~ojc;  //complement 
assign JAD =  AAD & EAB  |  ABD & EBB  |  ACD & ECB  |  ADD & EDB  ; 
assign jad = ~JAD;  //complement 
assign JED =  AAD & EAB  |  ABD & EBB  |  ACD & ECB  |  ADD & EDB  ; 
assign jed = ~JED; //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign rcd = ~RCD;  //complement 
assign rgd = ~RGD;  //complement 
assign LAD = ~lad;  //complement 
assign OJD = ~ojd;  //complement 
assign JBC =  AEC & EEB  |  AFC & EFB  |  AGC & EGB  |  AHC & EHB  ; 
assign jbc = ~JBC;  //complement 
assign JFC =  AEC & EEB  |  AFC & EFB  |  AGC & EGB  |  AHC & EHB  ; 
assign jfc = ~JFC; //complement 
assign afc = ~AFC;  //complement 
assign afd = ~AFD;  //complement 
assign ogc = ~OGC;  //complement 
assign oic = ~OIC;  //complement 
assign sac = ~SAC;  //complement 
assign oac = ~OAC;  //complement 
assign occ = ~OCC;  //complement 
assign oec = ~OEC;  //complement 
assign JBD =  AED & EEB  |  AFD & EFB  |  AGD & EGB  |  AHD & EHB  ; 
assign jbd = ~JBD;  //complement 
assign JFD =  AED & EEB  |  AFD & EFB  |  AGD & EGB  |  AHD & EHB  ; 
assign jfd = ~JFD; //complement 
assign ahc = ~AHC;  //complement 
assign ahd = ~AHD;  //complement 
assign ogd = ~OGD;  //complement 
assign oid = ~OID;  //complement 
assign sad = ~SAD;  //complement 
assign oad = ~OAD;  //complement 
assign ocd = ~OCD;  //complement 
assign oed = ~OED;  //complement 
assign JCC =  AIC & EIB  |  AJC & EJB  |  AKC & EKB  |  ALC & ELB  ; 
assign jcc = ~JCC;  //complement 
assign JGC =  AIC & EIB  |  AJC & EJB  |  AKC & EKB  |  ALC & ELB  ; 
assign jgc = ~JGC; //complement 
assign ajc = ~AJC;  //complement 
assign ajd = ~AJD;  //complement 
assign ohc = ~OHC;  //complement 
assign sbc = ~SBC;  //complement 
assign obc = ~OBC;  //complement 
assign odc = ~ODC;  //complement 
assign ofc = ~OFC;  //complement 
assign JCD =  AID & EIB  |  AJD & EJB  |  AKD & EKB  |  ALD & ELB  ; 
assign jcd = ~JCD;  //complement 
assign JGD =  AID & EIB  |  AJD & EJB  |  AKD & EKB  |  ALD & ELB  ; 
assign jgd = ~JGD; //complement 
assign alc = ~ALC;  //complement 
assign ald = ~ALD;  //complement 
assign ohd = ~OHD;  //complement 
assign sbd = ~SBD;  //complement 
assign obd = ~OBD;  //complement 
assign odd = ~ODD;  //complement 
assign ofd = ~OFD;  //complement 
assign JDC =  AMC & EMB  |  ANC & ENB  |  AOC & EOB  |  APC & EPB  ; 
assign jdc = ~JDC;  //complement 
assign JHC =  AMC & EMB  |  ANC & ENB  |  AOC & EOB  |  APC & EPB  ; 
assign jhc = ~JHC; //complement 
assign anc = ~ANC;  //complement 
assign and = ~AND;  //complement 
assign rdc = ~RDC;  //complement 
assign rhc = ~RHC;  //complement 
assign ome = ~OME;  //complement 
assign JDD =  AMD & EMB  |  AND & ENB  |  AOD & EOB  |  APD & EPB  ; 
assign jdd = ~JDD;  //complement 
assign JHD =  AMD & EMB  |  AND & ENB  |  AOD & EOB  |  APD & EPB  ; 
assign jhd = ~JHD; //complement 
assign apc = ~APC;  //complement 
assign apd = ~APD;  //complement 
assign rdd = ~RDD;  //complement 
assign rhd = ~RHD;  //complement 
assign omf = ~OMF;  //complement 
assign GBB =  CBA  ; 
assign gbb = ~GBB;  //complement 
assign GBC =  CBA & DBB  |  CBB  ; 
assign gbc = ~GBC;  //complement 
assign cba = ~CBA;  //complement 
assign dba = ~DBA;  //complement 
assign GBD =  CBA & DBB & DBC  |  CBB & DBC  |  CBC  ; 
assign gbd = ~GBD;  //complement 
assign cbb = ~CBB;  //complement 
assign dbb = ~DBB;  //complement 
assign KBA = ~kba;  //complement 
assign KBE = ~kbe;  //complement 
assign GBE =  CBA & DBB & DBC & DBD  |  CBB & DBC & DBD  |  CBC & DBD  |  CBD  ; 
assign gbe = ~GBE;  //complement 
assign KBB = ~kbb;  //complement 
assign KBF = ~kbf;  //complement 
assign MAB = ~mab;  //complement 
assign NAB = ~nab;  //complement 
assign KFB = ~kfb;  //complement 
assign KFF = ~kff;  //complement 
assign MAF = ~maf;  //complement 
assign NAF = ~naf;  //complement 
assign KFA = ~kfa;  //complement 
assign KFE = ~kfe;  //complement 
assign GFE =  CFA & DFB & DFC & DFD  |  CFB & DFC & DFD  |  CFC & DFD  |  CFD  ; 
assign gfe = ~GFE;  //complement 
assign omg = ~OMG;  //complement 
assign GFD =  CFA & DFB & DFC  |  CFB & DFC  |  CFC  ; 
assign gfd = ~GFD;  //complement 
assign cfa = ~CFA;  //complement 
assign dfa = ~DFA;  //complement 
assign omh = ~OMH;  //complement 
assign GFB =  CFA  ; 
assign gfb = ~GFB;  //complement 
assign GFC =  CFA & DFB  |  CFB  ; 
assign gfc = ~GFC;  //complement 
assign cfb = ~CFB;  //complement 
assign dfb = ~DFB;  //complement 
assign bba = ~BBA;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign bbb = ~BBB;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign eac = ~EAC;  //complement 
assign ebc = ~EBC;  //complement 
assign ecc = ~ECC;  //complement 
assign edc = ~EDC;  //complement 
assign rae = ~RAE;  //complement 
assign raf = ~RAF;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign jia =  saa & sab & sac & sad  ; 
assign JIA = ~jia;  //complement  
assign jib =  sae & saf & sag & sah  ; 
assign JIB = ~jib;  //complement 
assign REE = RAE; 
assign ree = ~REE; //complement 
assign REF = RAF; 
assign ref = ~REF;  //complement 
assign RIE = RAE; 
assign rie = ~RIE;  //complement 
assign RIF = RAF; 
assign rif = ~RIF;  //complement 
assign tab = ~TAB;  //complement 
assign taj = ~TAJ;  //complement 
assign tkb = ~TKB;  //complement 
assign tkj = ~TKJ;  //complement 
assign age = ~AGE;  //complement 
assign agf = ~AGF;  //complement 
assign eec = ~EEC;  //complement 
assign efc = ~EFC;  //complement 
assign egc = ~EGC;  //complement 
assign ehc = ~EHC;  //complement 
assign RFE = RBE; 
assign rfe = ~RFE; //complement 
assign RFF = RBF; 
assign rff = ~RFF;  //complement 
assign RJE = RBE; 
assign rje = ~RJE;  //complement 
assign RJF = RBF; 
assign rjf = ~RJF;  //complement 
assign taf = ~TAF;  //complement 
assign tan = ~TAN;  //complement 
assign tkf = ~TKF;  //complement 
assign tkn = ~TKN;  //complement 
assign aie = ~AIE;  //complement 
assign aif = ~AIF;  //complement 
assign EIC = ~eic;  //complement 
assign EJC = ~ejc;  //complement 
assign EKC = ~ekc;  //complement 
assign rbe = ~RBE;  //complement 
assign rbf = ~RBF;  //complement 
assign ake = ~AKE;  //complement 
assign akf = ~AKF;  //complement 
assign ELC = ~elc;  //complement 
assign EPC = ~epc;  //complement 
assign bfa = ~BFA;  //complement 
assign ame = ~AME;  //complement 
assign amf = ~AMF;  //complement 
assign EMC = ~emc;  //complement 
assign ENC = ~enc;  //complement 
assign EOC = ~eoc;  //complement 
assign bfb = ~BFB;  //complement 
assign aoe = ~AOE;  //complement 
assign aof = ~AOF;  //complement 
assign jie =  sba & sbb & sbc & sbd & scm & scn  ; 
assign JIE = ~jie;  //complement  
assign jif =  sbe & sbf & sbg & sbh  ; 
assign JIF = ~jif;  //complement 
assign JAE =  AAE & EAC  |  ABE & EBC  |  ACE & ECC  |  ADE & EDC  ; 
assign jae = ~JAE;  //complement 
assign JEE =  AAE & EAC  |  ABE & EBC  |  ACE & ECC  |  ADE & EDC  ; 
assign jee = ~JEE; //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign rce = ~RCE;  //complement 
assign rge = ~RGE;  //complement 
assign LAE = ~lae;  //complement 
assign OJE = ~oje;  //complement 
assign JAF =  AAF & EAC  |  ABF & EBC  |  ACF & ECC  |  ADF & EDC  ; 
assign jaf = ~JAF;  //complement 
assign JEF =  AAF & EAC  |  ABF & EBC  |  ACF & ECC  |  ADF & EDC  ; 
assign jef = ~JEF; //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign rcf = ~RCF;  //complement 
assign rgf = ~RGF;  //complement 
assign LAF = ~laf;  //complement 
assign OJF = ~ojf;  //complement 
assign JBE =  AEE & EEC  |  AFE & EFC  |  AGE & EGC  |  AHE & EHC  ; 
assign jbe = ~JBE;  //complement 
assign JFE =  AEE & EEC  |  AFE & EFC  |  AGE & EGC  |  AHE & EHC  ; 
assign jfe = ~JFE; //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign oge = ~OGE;  //complement 
assign oie = ~OIE;  //complement 
assign sae = ~SAE;  //complement 
assign oae = ~OAE;  //complement 
assign oce = ~OCE;  //complement 
assign oee = ~OEE;  //complement 
assign JBF =  AEF & EEC  |  AFF & EFC  |  AGF & EGC  |  AHF & EHC  ; 
assign jbf = ~JBF;  //complement 
assign JFF =  AEF & EEC  |  AFF & EFC  |  AGF & EGC  |  AHF & EHC  ; 
assign jff = ~JFF; //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign ogf = ~OGF;  //complement 
assign oif = ~OIF;  //complement 
assign saf = ~SAF;  //complement 
assign oaf = ~OAF;  //complement 
assign ocf = ~OCF;  //complement 
assign oef = ~OEF;  //complement 
assign JCE =  AIE & EIC  |  AJE & EJC  |  AKE & EKC  |  ALE & ELC  ; 
assign jce = ~JCE;  //complement 
assign JGE =  AIE & EIC  |  AJE & EJC  |  AKE & EKC  |  ALE & ELC  ; 
assign jge = ~JGE; //complement 
assign aje = ~AJE;  //complement 
assign ajf = ~AJF;  //complement 
assign ohe = ~OHE;  //complement 
assign sbe = ~SBE;  //complement 
assign obe = ~OBE;  //complement 
assign ode = ~ODE;  //complement 
assign ofe = ~OFE;  //complement 
assign JCF =  AIF & EIC  |  AJF & EJC  |  AKF & EKC  |  ALF & ELC  ; 
assign jcf = ~JCF;  //complement 
assign JGF =  AIF & EIC  |  AJF & EJC  |  AKF & EKC  |  ALF & ELC  ; 
assign jgf = ~JGF; //complement 
assign ale = ~ALE;  //complement 
assign alf = ~ALF;  //complement 
assign ohf = ~OHF;  //complement 
assign sbf = ~SBF;  //complement 
assign obf = ~OBF;  //complement 
assign odf = ~ODF;  //complement 
assign off = ~OFF;  //complement 
assign JDE =  AME & EMC  |  ANE & ENC  |  AOE & EOC  |  APE & EPC  ; 
assign jde = ~JDE;  //complement 
assign JHE =  AME & EMC  |  ANE & ENC  |  AOE & EOC  |  APE & EPC  ; 
assign jhe = ~JHE; //complement 
assign ane = ~ANE;  //complement 
assign anf = ~ANF;  //complement 
assign rde = ~RDE;  //complement 
assign rhe = ~RHE;  //complement 
assign tcg = qcc; 
assign TCG = ~tcg; //complement 
assign tch = qcc; 
assign TCH = ~tch;  //complement 
assign tdg = qcd; 
assign TDG = ~tdg;  //complement 
assign tdh = qcd; 
assign TDH = ~tdh;  //complement 
assign JDF =  AMF & EMC  |  ANF & ENC  |  AOF & EOC  |  APF & EPC  ; 
assign jdf = ~JDF;  //complement 
assign JHF =  AMF & EMC  |  ANF & ENC  |  AOF & EOC  |  APF & EPC  ; 
assign jhf = ~JHF; //complement 
assign ape = ~APE;  //complement 
assign apf = ~APF;  //complement 
assign rdf = ~RDF;  //complement 
assign rhf = ~RHF;  //complement 
assign teg = qce; 
assign TEG = ~teg; //complement 
assign teh = qce; 
assign TEH = ~teh;  //complement 
assign tfg = qcf; 
assign TFG = ~tfg;  //complement 
assign tfh = qcf; 
assign TFH = ~tfh;  //complement 
assign gbf =  dba  ; 
assign GBF = ~gbf;  //complement 
assign gbg =  dba & cbb  |  dbb  ; 
assign GBG = ~gbg;  //complement 
assign cbc = ~CBC;  //complement 
assign dbc = ~DBC;  //complement 
assign gbh =  dba & cbb & cbc  |  dbb & cbc  |  dbc  ; 
assign GBH = ~gbh;  //complement 
assign cbd = ~CBD;  //complement 
assign dbd = ~DBD;  //complement 
assign KBC = ~kbc;  //complement 
assign KBG = ~kbg;  //complement 
assign HBA =  DBA & cba  ; 
assign hba = ~HBA;  //complement 
assign HBB =  DBB & cbb  ; 
assign hbb = ~HBB;  //complement 
assign HBC =  DBC & cbc  ; 
assign hbc = ~HBC;  //complement 
assign PAB =  QAE & NAA  |  MAA  ; 
assign pab = ~PAB;  //complement 
assign KBD = ~kbd;  //complement 
assign KBH = ~kbh;  //complement 
assign HBD =  DBD & cbd  ; 
assign hbd = ~HBD;  //complement  
assign HBE =  DBA & DBB & DBC & DBD  ; 
assign hbe = ~HBE;  //complement 
assign tja = ~TJA;  //complement 
assign tjb = ~TJB;  //complement 
assign tjc = ~TJC;  //complement 
assign tjd = ~TJD;  //complement 
assign KFD = ~kfd;  //complement 
assign KFH = ~kfh;  //complement 
assign HFD =  DFD & cfd  ; 
assign hfd = ~HFD;  //complement  
assign HFE =  DFA & DFB & DFC & DFD  ; 
assign hfe = ~HFE;  //complement 
assign tje = ~TJE;  //complement 
assign tjf = ~TJF;  //complement 
assign tjg = ~TJG;  //complement 
assign tjh = ~TJH;  //complement 
assign KFC = ~kfc;  //complement 
assign KFG = ~kfg;  //complement 
assign HFA =  DFA & cfa  ; 
assign hfa = ~HFA;  //complement 
assign HFB =  DFB & cfb  ; 
assign hfb = ~HFB;  //complement 
assign HFC =  DFC & cfc  ; 
assign hfc = ~HFC;  //complement 
assign PAF =  QAF & NAE  |  MAE  ; 
assign paf = ~PAF;  //complement 
assign gfh =  dfa & cfb & cfc  |  dfb & cfc  |  dfc  ; 
assign GFH = ~gfh;  //complement 
assign cfc = ~CFC;  //complement 
assign dfc = ~DFC;  //complement 
assign gff =  dfa  ; 
assign GFF = ~gff;  //complement 
assign gfg =  dfa & cfb  |  dfb  ; 
assign GFG = ~gfg;  //complement 
assign cfd = ~CFD;  //complement 
assign dfd = ~DFD;  //complement 
assign bbc = ~BBC;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign QFE = ~qfe;  //complement 
assign QFF = ~qff;  //complement 
assign QFG = ~qfg;  //complement 
assign bbd = ~BBD;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign ead = ~EAD;  //complement 
assign ebd = ~EBD;  //complement 
assign ecd = ~ECD;  //complement 
assign edd = ~EDD;  //complement 
assign rag = ~RAG;  //complement 
assign rah = ~RAH;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign qfb = ~QFB;  //complement 
assign qfc = ~QFC;  //complement 
assign REG = RAG; 
assign reg = ~REG; //complement 
assign REH = RAH; 
assign reh = ~REH;  //complement 
assign RIG = RAG; 
assign rig = ~RIG;  //complement 
assign RIH = RAH; 
assign rih = ~RIH;  //complement 
assign taa = ~TAA;  //complement 
assign tai = ~TAI;  //complement 
assign tka = ~TKA;  //complement 
assign tki = ~TKI;  //complement 
assign agg = ~AGG;  //complement 
assign agh = ~AGH;  //complement 
assign eed = ~EED;  //complement 
assign efd = ~EFD;  //complement 
assign egd = ~EGD;  //complement 
assign ehd = ~EHD;  //complement 
assign RFG = RBG; 
assign rfg = ~RFG; //complement 
assign RFH = RBH; 
assign rfh = ~RFH;  //complement 
assign RJG = RBG; 
assign rjg = ~RJG;  //complement 
assign RJH = RBH; 
assign rjh = ~RJH;  //complement 
assign tae = ~TAE;  //complement 
assign tam = ~TAM;  //complement 
assign tke = ~TKE;  //complement 
assign tkm = ~TKM;  //complement 
assign aig = ~AIG;  //complement 
assign aih = ~AIH;  //complement 
assign EID = ~eid;  //complement 
assign EJD = ~ejd;  //complement 
assign EKD = ~ekd;  //complement 
assign rbg = ~RBG;  //complement 
assign rbh = ~RBH;  //complement 
assign akg = ~AKG;  //complement 
assign akh = ~AKH;  //complement 
assign ELD = ~eld;  //complement 
assign EPD = ~epd;  //complement 
assign bfc = ~BFC;  //complement 
assign amg = ~AMG;  //complement 
assign amh = ~AMH;  //complement 
assign EMD = ~emd;  //complement 
assign END = ~end;  //complement 
assign EOD = ~eod;  //complement 
assign bfd = ~BFD;  //complement 
assign aog = ~AOG;  //complement 
assign aoh = ~AOH;  //complement 
assign tbe = ~TBE;  //complement 
assign tbf = ~TBF;  //complement 
assign tbg = ~TBG;  //complement 
assign tbh = ~TBH;  //complement 
assign JAG =  AAG & EAD  |  ABG & EBD  |  ACG & ECD  |  ADG & EDD  ; 
assign jag = ~JAG;  //complement 
assign JEG =  AAG & EAD  |  ABG & EBD  |  ACG & ECD  |  ADG & EDD  ; 
assign jeg = ~JEG; //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign rcg = ~RCG;  //complement 
assign rgg = ~RGG;  //complement 
assign TCE = QCC; 
assign tce = ~TCE; //complement 
assign TCF = QCC; 
assign tcf = ~TCF;  //complement 
assign TDE = QCD; 
assign tde = ~TDE;  //complement 
assign TDF = QCD; 
assign tdf = ~TDF;  //complement 
assign JAH =  AAH & EAD  |  ABH & EBD  |  ACH & ECD  |  ADH & EDD  ; 
assign jah = ~JAH;  //complement 
assign JEH =  AAH & EAD  |  ABH & EBD  |  ACH & ECD  |  ADH & EDD  ; 
assign jeh = ~JEH; //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign rch = ~RCH;  //complement 
assign rgh = ~RGH;  //complement 
assign TEE = QCE; 
assign tee = ~TEE; //complement 
assign TEF = QCE; 
assign tef = ~TEF;  //complement 
assign TFE = QCF; 
assign tfe = ~TFE;  //complement 
assign TFF = QCF; 
assign tff = ~TFF;  //complement 
assign JBG =  AEG & EED  |  AFG & EFD  |  AGG & EGD  |  AHG & EHD  ; 
assign jbg = ~JBG;  //complement 
assign JFG =  AEG & EED  |  AFG & EFD  |  AGG & EGD  |  AHG & EHD  ; 
assign jfg = ~JFG; //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign ogg = ~OGG;  //complement 
assign oig = ~OIG;  //complement 
assign sag = ~SAG;  //complement 
assign oag = ~OAG;  //complement 
assign ocg = ~OCG;  //complement 
assign oeg = ~OEG;  //complement 
assign JBH =  AEH & EED  |  AFH & EFD  |  AGH & EGD  |  AHH & EHD  ; 
assign jbh = ~JBH;  //complement 
assign JFH =  AEH & EED  |  AFH & EFD  |  AGH & EGD  |  AHH & EHD  ; 
assign jfh = ~JFH; //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign ogh = ~OGH;  //complement 
assign oih = ~OIH;  //complement 
assign sah = ~SAH;  //complement 
assign oah = ~OAH;  //complement 
assign och = ~OCH;  //complement 
assign oeh = ~OEH;  //complement 
assign JCG =  AIG & EID  |  AJG & EJD  |  AKG & EKD  |  ALG & ELD  ; 
assign jcg = ~JCG;  //complement 
assign JGG =  AIG & EID  |  AJG & EJD  |  AKG & EKD  |  ALG & ELD  ; 
assign jgg = ~JGG; //complement 
assign ajg = ~AJG;  //complement 
assign ajh = ~AJH;  //complement 
assign ohg = ~OHG;  //complement 
assign sbg = ~SBG;  //complement 
assign obg = ~OBG;  //complement 
assign odg = ~ODG;  //complement 
assign ofg = ~OFG;  //complement 
assign JCH =  AIH & EID  |  AJH & EJD  |  AKH & EKD  |  ALH & ELD  ; 
assign jch = ~JCH;  //complement 
assign JGH =  AIH & EID  |  AJH & EJD  |  AKH & EKD  |  ALH & ELD  ; 
assign jgh = ~JGH; //complement 
assign alg = ~ALG;  //complement 
assign alh = ~ALH;  //complement 
assign ohh = ~OHH;  //complement 
assign sbh = ~SBH;  //complement 
assign obh = ~OBH;  //complement 
assign odh = ~ODH;  //complement 
assign ofh = ~OFH;  //complement 
assign JDG =  AMG & EMD  |  ANG & END  |  AOG & EOD  |  APG & EPD  ; 
assign jdg = ~JDG;  //complement 
assign JHG =  AMG & EMD  |  ANG & END  |  AOG & EOD  |  APG & EPD  ; 
assign jhg = ~JHG; //complement 
assign ang = ~ANG;  //complement 
assign anh = ~ANH;  //complement 
assign rdg = ~RDG;  //complement 
assign rhg = ~RHG;  //complement 
assign FAA = ~QDC & ~QDB & ~QDA  ; 
assign FAB = ~QDC & ~QDB &  QDA  ; 
assign FAC = ~QDC &  QDB & ~QDA  ; 
assign FAD = ~QDC &  QDB &  QDA  ; 
assign FAE =  QDC & ~QDB & ~QDA  ; 
assign FAF =  QDC & ~QDB &  QDA ; 
assign FAG =  QDC &  QDB & ~QDA  ; 
assign FAH =  QDC &  QDB &  QDA ; 
assign FAI = ZZI ; 
assign JDH =  AMH & EMD  |  ANH & END  |  AOH & EOD  |  APH & EPD  ; 
assign jdh = ~JDH;  //complement 
assign JHH =  AMH & EMD  |  ANH & END  |  AOH & EOD  |  APH & EPD  ; 
assign jhh = ~JHH; //complement 
assign apg = ~APG;  //complement 
assign aph = ~APH;  //complement 
assign rdh = ~RDH;  //complement 
assign rhh = ~RHH;  //complement 
assign FBA = ~QDC & ~QDB & ~QDA  ; 
assign FBB = ~QDC & ~QDB &  QDA  ; 
assign FBC = ~QDC &  QDB & ~QDA  ; 
assign FBD = ~QDC &  QDB &  QDA  ; 
assign FBE =  QDC & ~QDB & ~QDA  ; 
assign FBF =  QDC & ~QDB &  QDA ; 
assign FBG =  QDC &  QDB & ~QDA  ; 
assign FBH =  QDC &  QDB &  QDA ; 
assign FBI = ZZI ; 
assign GCB =  CCA  ; 
assign gcb = ~GCB;  //complement 
assign GCC =  CCA & DCB  |  CCB  ; 
assign gcc = ~GCC;  //complement 
assign cca = ~CCA;  //complement 
assign dca = ~DCA;  //complement 
assign GCD =  CCA & DCB & DCC  |  CCB & DCC  |  CCC  ; 
assign gcd = ~GCD;  //complement 
assign ccb = ~CCB;  //complement 
assign dcb = ~DCB;  //complement 
assign KCA = ~kca;  //complement 
assign KCE = ~kce;  //complement 
assign GCE =  CCA & DCB & DCC & DCD  |  CCB & DCC & DCD  |  CCC & DCD  |  CCD  ; 
assign gce = ~GCE;  //complement 
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign tic = ~TIC;  //complement 
assign tid = ~TID;  //complement 
assign KCB = ~kcb;  //complement 
assign KCF = ~kcf;  //complement 
assign MAC = ~mac;  //complement 
assign NAC = ~nac;  //complement 
assign KGB = ~kgb;  //complement 
assign KGF = ~kgf;  //complement 
assign MAG = ~mag;  //complement 
assign NAG = ~nag;  //complement 
assign KGA = ~kga;  //complement 
assign KGE = ~kge;  //complement 
assign GGE =  CGA & DGB & DGC & DGD  |  CGB & DGC & DGD  |  CGC & DGD  |  CGD  ; 
assign gge = ~GGE;  //complement 
assign tie = ~TIE;  //complement 
assign tif = ~TIF;  //complement 
assign tig = ~TIG;  //complement 
assign tih = ~TIH;  //complement 
assign GGD =  CGA & DGB & DGC  |  CGB & DGC  |  CGC  ; 
assign ggd = ~GGD;  //complement 
assign cga = ~CGA;  //complement 
assign dga = ~DGA;  //complement 
assign GGB =  CGA  ; 
assign ggb = ~GGB;  //complement 
assign GGC =  CGA & DGB  |  CGB  ; 
assign ggc = ~GGC;  //complement 
assign cgb = ~CGB;  //complement 
assign dgb = ~DGB;  //complement 
assign bca = ~BCA;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign QHA = QEA; 
assign qha = ~QHA; //complement 
assign QHB = QEB; 
assign qhb = ~QHB;  //complement 
assign QIA = QEA; 
assign qia = ~QIA;  //complement 
assign QIB = QEB; 
assign qib = ~QIB;  //complement 
assign bcb = ~BCB;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign eae = ~EAE;  //complement 
assign ebe = ~EBE;  //complement 
assign ece = ~ECE;  //complement 
assign ede = ~EDE;  //complement 
assign rai = ~RAI;  //complement 
assign raj = ~RAJ;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign REI = RAI; 
assign rei = ~REI; //complement 
assign REJ = RAJ; 
assign rej = ~REJ;  //complement 
assign RII = RAI; 
assign rii = ~RII;  //complement 
assign RIJ = RAJ; 
assign rij = ~RIJ;  //complement 
assign tla = ~TLA;  //complement 
assign tli = ~TLI;  //complement 
assign tma = ~TMA;  //complement 
assign tmi = ~TMI;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign eee = ~EEE;  //complement 
assign efe = ~EFE;  //complement 
assign ege = ~EGE;  //complement 
assign ehe = ~EHE;  //complement 
assign RFI = RBI; 
assign rfi = ~RFI; //complement 
assign RFJ = RBJ; 
assign rfj = ~RFJ;  //complement 
assign RJI = RBI; 
assign rji = ~RJI;  //complement 
assign RJJ = RBJ; 
assign rjj = ~RJJ;  //complement 
assign tle = ~TLE;  //complement 
assign tlm = ~TLM;  //complement 
assign tme = ~TME;  //complement 
assign tmm = ~TMM;  //complement 
assign aii = ~AII;  //complement 
assign aij = ~AIJ;  //complement 
assign EIE = ~eie;  //complement 
assign EJE = ~eje;  //complement 
assign EKE = ~eke;  //complement 
assign rbi = ~RBI;  //complement 
assign rbj = ~RBJ;  //complement 
assign aki = ~AKI;  //complement 
assign akj = ~AKJ;  //complement 
assign ELE = ~ele;  //complement 
assign EPE = ~epe;  //complement 
assign bga = ~BGA;  //complement 
assign ami = ~AMI;  //complement 
assign amj = ~AMJ;  //complement 
assign EME = ~eme;  //complement 
assign ENE = ~ene;  //complement 
assign EOE = ~eoe;  //complement 
assign bgb = ~BGB;  //complement 
assign aoi = ~AOI;  //complement 
assign aoj = ~AOJ;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tbc = ~TBC;  //complement 
assign tbd = ~TBD;  //complement 
assign JAI =  AAI & EAE  |  ABI & EBE  |  ACI & ECE  |  ADI & EDE  ; 
assign jai = ~JAI;  //complement 
assign JEI =  AAI & EAE  |  ABI & EBE  |  ACI & ECE  |  ADI & EDE  ; 
assign jei = ~JEI; //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign rci = ~RCI;  //complement 
assign rgi = ~RGI;  //complement 
assign QEA = ~qea;  //complement 
assign QEB = ~qeb;  //complement 
assign JAJ =  AAJ & EAE  |  ABJ & EBE  |  ACJ & ECE  |  ADJ & EDE  ; 
assign jaj = ~JAJ;  //complement 
assign JEJ =  AAJ & EAE  |  ABJ & EBE  |  ACJ & ECE  |  ADJ & EDE  ; 
assign jej = ~JEJ; //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign rcj = ~RCJ;  //complement 
assign rgj = ~RGJ;  //complement 
assign qaa = ~QAA;  //complement 
assign qfa = ~QFA;  //complement 
assign qfh = ~QFH;  //complement 
assign JBI =  AEI & EEE  |  AFI & EFE  |  AGI & EGE  |  AHI & EHE  ; 
assign jbi = ~JBI;  //complement 
assign JFI =  AEI & EEE  |  AFI & EFE  |  AGI & EGE  |  AHI & EHE  ; 
assign jfi = ~JFI; //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign ogi = ~OGI;  //complement 
assign sai = ~SAI;  //complement 
assign oai = ~OAI;  //complement 
assign oci = ~OCI;  //complement 
assign oei = ~OEI;  //complement 
assign JBJ =  AEJ & EEE  |  AFJ & EFE  |  AGJ & EGE  |  AHJ & EHE  ; 
assign jbj = ~JBJ;  //complement 
assign JFJ =  AEJ & EEE  |  AFJ & EFE  |  AGJ & EGE  |  AHJ & EHE  ; 
assign jfj = ~JFJ; //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign ogj = ~OGJ;  //complement 
assign saj = ~SAJ;  //complement 
assign oaj = ~OAJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign oej = ~OEJ;  //complement 
assign JCI =  AII & EIE  |  AJI & EJE  |  AKI & EKE  |  ALI & ELE  ; 
assign jci = ~JCI;  //complement 
assign JGI =  AII & EIE  |  AJI & EJE  |  AKI & EKE  |  ALI & ELE  ; 
assign jgi = ~JGI; //complement 
assign aji = ~AJI;  //complement 
assign ajj = ~AJJ;  //complement 
assign ohi = ~OHI;  //complement 
assign sbi = ~SBI;  //complement 
assign obi = ~OBI;  //complement 
assign odi = ~ODI;  //complement 
assign ofi = ~OFI;  //complement 
assign JCJ =  AIJ & EIE  |  AJJ & EJE  |  AKJ & EKE  |  ALJ & ELE  ; 
assign jcj = ~JCJ;  //complement 
assign JGJ =  AIJ & EIE  |  AJJ & EJE  |  AKJ & EKE  |  ALJ & ELE  ; 
assign jgj = ~JGJ; //complement 
assign ali = ~ALI;  //complement 
assign alj = ~ALJ;  //complement 
assign ohj = ~OHJ;  //complement 
assign sbj = ~SBJ;  //complement 
assign obj = ~OBJ;  //complement 
assign odj = ~ODJ;  //complement 
assign ofj = ~OFJ;  //complement 
assign JDI =  AMI & EME  |  ANI & ENE  |  AOI & EOE  |  API & EPE  ; 
assign jdi = ~JDI;  //complement 
assign JHI =  AMI & EME  |  ANI & ENE  |  AOI & EOE  |  API & EPE  ; 
assign jhi = ~JHI; //complement 
assign ani = ~ANI;  //complement 
assign anj = ~ANJ;  //complement 
assign rdi = ~RDI;  //complement 
assign rhi = ~RHI;  //complement 
assign QCA = ~qca;  //complement 
assign QCB = ~qcb;  //complement 
assign JDJ =  AMJ & EME  |  ANJ & ENE  |  AOJ & EOE  |  APJ & EPE  ; 
assign jdj = ~JDJ;  //complement 
assign JHJ =  AMJ & EME  |  ANJ & ENE  |  AOJ & EOE  |  APJ & EPE  ; 
assign jhj = ~JHJ; //complement 
assign api = ~API;  //complement 
assign apj = ~APJ;  //complement 
assign rdj = ~RDJ;  //complement 
assign rhj = ~RHJ;  //complement 
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign gcf =  dca  ; 
assign GCF = ~gcf;  //complement 
assign gcg =  dca & ccb  |  dcb  ; 
assign GCG = ~gcg;  //complement 
assign ccc = ~CCC;  //complement 
assign dcc = ~DCC;  //complement 
assign gch =  dca & ccb & ccc  |  dcb & ccc  |  dcc  ; 
assign GCH = ~gch;  //complement 
assign ccd = ~CCD;  //complement 
assign dcd = ~DCD;  //complement 
assign KCC = ~kcc;  //complement 
assign KCG = ~kcg;  //complement 
assign HCA =  DCA & cca  ; 
assign hca = ~HCA;  //complement 
assign HCB =  DCB & ccb  ; 
assign hcb = ~HCB;  //complement 
assign HCC =  DCC & ccc  ; 
assign hcc = ~HCC;  //complement 
assign PAC =  QAE & NAA & NAB  |  MAA & NAB  |  MAB  ; 
assign pac = ~PAC;  //complement 
assign KCD = ~kcd;  //complement 
assign KCH = ~kch;  //complement 
assign HCD =  DCD & ccd  ; 
assign hcd = ~HCD;  //complement  
assign HCE =  DCA & DCB & DCC & DCD  ; 
assign hce = ~HCE;  //complement 
assign KGD = ~kgd;  //complement 
assign KGH = ~kgh;  //complement 
assign HGD =  DGD & cgd  ; 
assign hgd = ~HGD;  //complement  
assign HGE =  DGA & DGB & DGC & DGD  ; 
assign hge = ~HGE;  //complement 
assign KGC = ~kgc;  //complement 
assign KGG = ~kgg;  //complement 
assign HGA =  DGA & cga  ; 
assign hga = ~HGA;  //complement 
assign HGB =  DGB & cgb  ; 
assign hgb = ~HGB;  //complement 
assign HGC =  DGC & cgc  ; 
assign hgc = ~HGC;  //complement 
assign PAG =  QAF & NAE & NAF  |  MAE & NAF  |  MAF  ; 
assign pag = ~PAG;  //complement 
assign ggh =  dga & cgb & cgc  |  dgb & cgc  |  dgc  ; 
assign GGH = ~ggh;  //complement 
assign cgc = ~CGC;  //complement 
assign dgc = ~DGC;  //complement 
assign ggf =  dga  ; 
assign GGF = ~ggf;  //complement 
assign ggg =  dga & cgb  |  dgb  ; 
assign GGG = ~ggg;  //complement 
assign cgd = ~CGD;  //complement 
assign dgd = ~DGD;  //complement 
assign bcc = ~BCC;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign QHC = QEC; 
assign qhc = ~QHC; //complement 
assign QHD = QED; 
assign qhd = ~QHD;  //complement 
assign QIC = QEC; 
assign qic = ~QIC;  //complement 
assign QID = QED; 
assign qid = ~QID;  //complement 
assign bcd = ~BCD;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign eaf = ~EAF;  //complement 
assign ebf = ~EBF;  //complement 
assign ecf = ~ECF;  //complement 
assign edf = ~EDF;  //complement 
assign rak = ~RAK;  //complement 
assign ral = ~RAL;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign qba = ~QBA;  //complement 
assign qbb = ~QBB;  //complement 
assign qbc = ~QBC;  //complement 
assign REK = RAK; 
assign rek = ~REK; //complement 
assign REL = RAL; 
assign rel = ~REL;  //complement 
assign RIK = RAK; 
assign rik = ~RIK;  //complement 
assign RIL = RAL; 
assign ril = ~RIL;  //complement 
assign tlb = ~TLB;  //complement 
assign tlj = ~TLJ;  //complement 
assign tmb = ~TMB;  //complement 
assign tmj = ~TMJ;  //complement 
assign agk = ~AGK;  //complement 
assign agl = ~AGL;  //complement 
assign eef = ~EEF;  //complement 
assign eff = ~EFF;  //complement 
assign egf = ~EGF;  //complement 
assign ehf = ~EHF;  //complement 
assign RFK = RBK; 
assign rfk = ~RFK; //complement 
assign RFL = RBL; 
assign rfl = ~RFL;  //complement 
assign RJK = RBK; 
assign rjk = ~RJK;  //complement 
assign RJL = RBL; 
assign rjl = ~RJL;  //complement 
assign tlf = ~TLF;  //complement 
assign tln = ~TLN;  //complement 
assign tmf = ~TMF;  //complement 
assign tmn = ~TMN;  //complement 
assign aik = ~AIK;  //complement 
assign ail = ~AIL;  //complement 
assign EIF = ~eif;  //complement 
assign EJF = ~ejf;  //complement 
assign EKF = ~ekf;  //complement 
assign rbk = ~RBK;  //complement 
assign rbl = ~RBL;  //complement 
assign akk = ~AKK;  //complement 
assign akl = ~AKL;  //complement 
assign ELF = ~elf;  //complement 
assign EPF = ~epf;  //complement 
assign bgc = ~BGC;  //complement 
assign amk = ~AMK;  //complement 
assign aml = ~AML;  //complement 
assign EMF = ~emf;  //complement 
assign ENF = ~enf;  //complement 
assign EOF = ~eof;  //complement 
assign bgd = ~BGD;  //complement 
assign aok = ~AOK;  //complement 
assign aol = ~AOL;  //complement 
assign JAK =  AAK & EAF  |  ABK & EBF  |  ACK & ECF  |  ADK & EDF  ; 
assign jak = ~JAK;  //complement 
assign JEK =  AAK & EAF  |  ABK & EBF  |  ACK & ECF  |  ADK & EDF  ; 
assign jek = ~JEK; //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign rck = ~RCK;  //complement 
assign rgk = ~RGK;  //complement 
assign QEC = ~qec;  //complement 
assign QED = ~qed;  //complement 
assign JAL =  AAL & EAF  |  ABL & EBF  |  ACL & ECF  |  ADL & EDF  ; 
assign jal = ~JAL;  //complement 
assign JEL =  AAL & EAF  |  ABL & EBF  |  ACL & ECF  |  ADL & EDF  ; 
assign jel = ~JEL; //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign rcl = ~RCL;  //complement 
assign rgl = ~RGL;  //complement 
assign TCA = QCC; 
assign tca = ~TCA; //complement 
assign TCB = QCC; 
assign tcb = ~TCB;  //complement 
assign TDA = QCD; 
assign tda = ~TDA;  //complement 
assign TDB = QCD; 
assign tdb = ~TDB;  //complement 
assign JBK =  AEK & EEF  |  AFK & EFF  |  AGK & EGF  |  AHK & EHF  ; 
assign jbk = ~JBK;  //complement 
assign JFK =  AEK & EEF  |  AFK & EFF  |  AGK & EGF  |  AHK & EHF  ; 
assign jfk = ~JFK; //complement 
assign afk = ~AFK;  //complement 
assign afl = ~AFL;  //complement 
assign ogk = ~OGK;  //complement 
assign sak = ~SAK;  //complement 
assign oak = ~OAK;  //complement 
assign ock = ~OCK;  //complement 
assign oek = ~OEK;  //complement 
assign JBL =  AEL & EEF  |  AFL & EFF  |  AGL & EGF  |  AHL & EHF  ; 
assign jbl = ~JBL;  //complement 
assign JFL =  AEL & EEF  |  AFL & EFF  |  AGL & EGF  |  AHL & EHF  ; 
assign jfl = ~JFL; //complement 
assign ahk = ~AHK;  //complement 
assign ahl = ~AHL;  //complement 
assign ogl = ~OGL;  //complement 
assign sal = ~SAL;  //complement 
assign oal = ~OAL;  //complement 
assign ocl = ~OCL;  //complement 
assign oel = ~OEL;  //complement 
assign JCK =  AIK & EIF  |  AJK & EJF  |  AKK & EKF  |  ALK & ELF  ; 
assign jck = ~JCK;  //complement 
assign JGK =  AIK & EIF  |  AJK & EJF  |  AKK & EKF  |  ALK & ELF  ; 
assign jgk = ~JGK; //complement 
assign ajk = ~AJK;  //complement 
assign ajl = ~AJL;  //complement 
assign ohk = ~OHK;  //complement 
assign sbk = ~SBK;  //complement 
assign obk = ~OBK;  //complement 
assign odk = ~ODK;  //complement 
assign ofk = ~OFK;  //complement 
assign JCL =  AIL & EIF  |  AJL & EJF  |  AKL & EKF  |  ALL & ELF  ; 
assign jcl = ~JCL;  //complement 
assign JGL =  AIL & EIF  |  AJL & EJF  |  AKL & EKF  |  ALL & ELF  ; 
assign jgl = ~JGL; //complement 
assign alk = ~ALK;  //complement 
assign all = ~ALL;  //complement 
assign ohl = ~OHL;  //complement 
assign sbl = ~SBL;  //complement 
assign obl = ~OBL;  //complement 
assign odl = ~ODL;  //complement 
assign ofl = ~OFL;  //complement 
assign JDK =  AMK & EMF  |  ANK & ENF  |  AOK & EOF  |  APK & EPF  ; 
assign jdk = ~JDK;  //complement 
assign JHK =  AMK & EMF  |  ANK & ENF  |  AOK & EOF  |  APK & EPF  ; 
assign jhk = ~JHK; //complement 
assign ank = ~ANK;  //complement 
assign anl = ~ANL;  //complement 
assign rdk = ~RDK;  //complement 
assign rhk = ~RHK;  //complement 
assign QCC = ~qcc;  //complement 
assign QCD = ~qcd;  //complement 
assign JDL =  AML & EMF  |  ANL & ENF  |  AOL & EOF  |  APL & EPF  ; 
assign jdl = ~JDL;  //complement 
assign JHL =  AML & EMF  |  ANL & ENF  |  AOL & EOF  |  APL & EPF  ; 
assign jhl = ~JHL; //complement 
assign apk = ~APK;  //complement 
assign apl = ~APL;  //complement 
assign rdl = ~RDL;  //complement 
assign rhl = ~RHL;  //complement 
assign tcc = qcc; 
assign TCC = ~tcc; //complement 
assign tcd = qcc; 
assign TCD = ~tcd;  //complement 
assign tdc = qcd; 
assign TDC = ~tdc;  //complement 
assign tdd = qcd; 
assign TDD = ~tdd;  //complement 
assign GDB =  CDA  ; 
assign gdb = ~GDB;  //complement 
assign GDC =  CDA & DDB  |  CDB  ; 
assign gdc = ~GDC;  //complement 
assign cda = ~CDA;  //complement 
assign dda = ~DDA;  //complement 
assign GDD =  CDA & DDB & DDC  |  CDB & DDC  |  CDC  ; 
assign gdd = ~GDD;  //complement 
assign cdb = ~CDB;  //complement 
assign ddb = ~DDB;  //complement 
assign KDA = ~kda;  //complement 
assign KDE = ~kde;  //complement 
assign GDE =  CDA & DDB & DDC & DDD  |  CDB & DDC & DDD  |  CDC & DDD  |  CDD  ; 
assign gde = ~GDE;  //complement 
assign KDB = ~kdb;  //complement 
assign KDF = ~kdf;  //complement 
assign qae = ~QAE;  //complement 
assign KHB = ~khb;  //complement 
assign KHF = ~khf;  //complement 
assign qaf = ~QAF;  //complement 
assign KHA = ~kha;  //complement 
assign KHE = ~khe;  //complement 
assign GHD =  CHA & DHB & DHC  |  CHB & DHC  |  CHC  ; 
assign ghd = ~GHD;  //complement 
assign cha = ~CHA;  //complement 
assign dha = ~DHA;  //complement 
assign GHB =  CHA  ; 
assign ghb = ~GHB;  //complement 
assign GHC =  CHA & DHB  |  CHB  ; 
assign ghc = ~GHC;  //complement 
assign chb = ~CHB;  //complement 
assign dhb = ~DHB;  //complement 
assign bda = ~BDA;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign QHE = QEE; 
assign qhe = ~QHE; //complement 
assign QHF = QEF; 
assign qhf = ~QHF;  //complement 
assign QIE = QEE; 
assign qie = ~QIE;  //complement 
assign QIF = QEF; 
assign qif = ~QIF;  //complement 
assign bdb = ~BDB;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign eag = ~EAG;  //complement 
assign ebg = ~EBG;  //complement 
assign ecg = ~ECG;  //complement 
assign edg = ~EDG;  //complement 
assign ram = ~RAM;  //complement 
assign ran = ~RAN;  //complement 
assign aem = ~AEM;  //complement 
assign aen = ~AEN;  //complement 
assign REM = RAM; 
assign rem = ~REM; //complement 
assign REN = RAN; 
assign ren = ~REN;  //complement 
assign RIM = RAM; 
assign rim = ~RIM;  //complement 
assign RIN = RAN; 
assign rin = ~RIN;  //complement 
assign tlc = ~TLC;  //complement 
assign tlk = ~TLK;  //complement 
assign tmc = ~TMC;  //complement 
assign tmk = ~TMK;  //complement 
assign agm = ~AGM;  //complement 
assign agn = ~AGN;  //complement 
assign eeg = ~EEG;  //complement 
assign efg = ~EFG;  //complement 
assign egg = ~EGG;  //complement 
assign ehg = ~EHG;  //complement 
assign RFM = RBM; 
assign rfm = ~RFM; //complement 
assign RFN = RBN; 
assign rfn = ~RFN;  //complement 
assign RJM = RBM; 
assign rjm = ~RJM;  //complement 
assign RJN = RBN; 
assign rjn = ~RJN;  //complement 
assign tlg = ~TLG;  //complement 
assign tlo = ~TLO;  //complement 
assign tmg = ~TMG;  //complement 
assign tmo = ~TMO;  //complement 
assign aim = ~AIM;  //complement 
assign ain = ~AIN;  //complement 
assign EIG = ~eig;  //complement 
assign EJG = ~ejg;  //complement 
assign EKG = ~ekg;  //complement 
assign rbm = ~RBM;  //complement 
assign rbn = ~RBN;  //complement 
assign akm = ~AKM;  //complement 
assign akn = ~AKN;  //complement 
assign ELG = ~elg;  //complement 
assign EPG = ~epg;  //complement 
assign bha = ~BHA;  //complement 
assign amm = ~AMM;  //complement 
assign amn = ~AMN;  //complement 
assign EMG = ~emg;  //complement 
assign ENG = ~eng;  //complement 
assign EOG = ~eog;  //complement 
assign bhb = ~BHB;  //complement 
assign aom = ~AOM;  //complement 
assign aon = ~AON;  //complement 
assign JAM =  AAM & EAG  |  ABM & EBG  |  ACM & ECG  |  ADM & EDG  ; 
assign jam = ~JAM;  //complement 
assign JEM =  AAM & EAG  |  ABM & EBG  |  ACM & ECG  |  ADM & EDG  ; 
assign jem = ~JEM; //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign rcm = ~RCM;  //complement 
assign rgm = ~RGM;  //complement 
assign QEE = ~qee;  //complement 
assign QEF = ~qef;  //complement 
assign JAN =  AAN & EAG  |  ABN & EBG  |  ACN & ECG  |  ADN & EDG  ; 
assign jan = ~JAN;  //complement 
assign JEN =  AAN & EAG  |  ABN & EBG  |  ACN & ECG  |  ADN & EDG  ; 
assign jen = ~JEN; //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign rcn = ~RCN;  //complement 
assign rgn = ~RGN;  //complement 
assign TEA = QCE; 
assign tea = ~TEA; //complement 
assign TEB = QCE; 
assign teb = ~TEB;  //complement 
assign TFA = QCF; 
assign tfa = ~TFA;  //complement 
assign TFB = QCF; 
assign tfb = ~TFB;  //complement 
assign JBM =  AEM & EEG  |  AFM & EFG  |  AGM & EGG  |  AHM & EHG  ; 
assign jbm = ~JBM;  //complement 
assign JFM =  AEM & EEG  |  AFM & EFG  |  AGM & EGG  |  AHM & EHG  ; 
assign jfm = ~JFM; //complement 
assign afm = ~AFM;  //complement 
assign afn = ~AFN;  //complement 
assign ogm = ~OGM;  //complement 
assign sam = ~SAM;  //complement 
assign oam = ~OAM;  //complement 
assign ocm = ~OCM;  //complement 
assign oem = ~OEM;  //complement 
assign JBN =  AEN & EEG  |  AFN & EFG  |  AGN & EGG  |  AHN & EHG  ; 
assign jbn = ~JBN;  //complement 
assign JFN =  AEN & EEG  |  AFN & EFG  |  AGN & EGG  |  AHN & EHG  ; 
assign jfn = ~JFN; //complement 
assign ahm = ~AHM;  //complement 
assign ahn = ~AHN;  //complement 
assign ogn = ~OGN;  //complement 
assign san = ~SAN;  //complement 
assign oan = ~OAN;  //complement 
assign ocn = ~OCN;  //complement 
assign oen = ~OEN;  //complement 
assign JCM =  AIM & EIG  |  AJM & EJG  |  AKM & EKG  |  ALM & ELG  ; 
assign jcm = ~JCM;  //complement 
assign JGM =  AIM & EIG  |  AJM & EJG  |  AKM & EKG  |  ALM & ELG  ; 
assign jgm = ~JGM; //complement 
assign ajm = ~AJM;  //complement 
assign ajn = ~AJN;  //complement 
assign ohm = ~OHM;  //complement 
assign sbm = ~SBM;  //complement 
assign scm = ~SCM;  //complement 
assign obm = ~OBM;  //complement 
assign odm = ~ODM;  //complement 
assign ofm = ~OFM;  //complement 
assign JCN =  AIN & EIG  |  AJN & EJG  |  AKN & EKG  |  ALN & ELG  ; 
assign jcn = ~JCN;  //complement 
assign JGN =  AIN & EIG  |  AJN & EJG  |  AKN & EKG  |  ALN & ELG  ; 
assign jgn = ~JGN; //complement 
assign alm = ~ALM;  //complement 
assign aln = ~ALN;  //complement 
assign ohn = ~OHN;  //complement 
assign sbn = ~SBN;  //complement 
assign scn = ~SCN;  //complement 
assign obn = ~OBN;  //complement 
assign odn = ~ODN;  //complement 
assign ofn = ~OFN;  //complement 
assign JDM =  AMM & EMG  |  ANM & ENG  |  AOM & EOG  |  APM & EPG  ; 
assign jdm = ~JDM;  //complement 
assign JHM =  AMM & EMG  |  ANM & ENG  |  AOM & EOG  |  APM & EPG  ; 
assign jhm = ~JHM; //complement 
assign anm = ~ANM;  //complement 
assign ann = ~ANN;  //complement 
assign rdm = ~RDM;  //complement 
assign rhm = ~RHM;  //complement 
assign QCE = ~qce;  //complement 
assign QCF = ~qcf;  //complement 
assign JDN =  AMN & EMG  |  ANN & ENG  |  AON & EOG  |  APN & EPG  ; 
assign jdn = ~JDN;  //complement 
assign JHN =  AMN & EMG  |  ANN & ENG  |  AON & EOG  |  APN & EPG  ; 
assign jhn = ~JHN; //complement 
assign apm = ~APM;  //complement 
assign apn = ~APN;  //complement 
assign rdn = ~RDN;  //complement 
assign rhn = ~RHN;  //complement 
assign tec = qce; 
assign TEC = ~tec; //complement 
assign ted = qce; 
assign TED = ~ted;  //complement 
assign tfc = qcf; 
assign TFC = ~tfc;  //complement 
assign tfd = qcf; 
assign TFD = ~tfd;  //complement 
assign gdf =  dda  ; 
assign GDF = ~gdf;  //complement 
assign gdg =  dda & cdb  |  ddb  ; 
assign GDG = ~gdg;  //complement 
assign cdc = ~CDC;  //complement 
assign ddc = ~DDC;  //complement 
assign gdh =  dda & cdb & cdc  |  ddb & cdc  |  ddc  ; 
assign GDH = ~gdh;  //complement 
assign cdd = ~CDD;  //complement 
assign ddd = ~DDD;  //complement 
assign KDC = ~kdc;  //complement 
assign KDG = ~kdg;  //complement 
assign HDA =  DDA & cda  ; 
assign hda = ~HDA;  //complement 
assign HDB =  DDB & cdb  ; 
assign hdb = ~HDB;  //complement 
assign HDC =  DDC & cdc  ; 
assign hdc = ~HDC;  //complement 
assign PAD =  QAE & NAA & NAB & NAC  |  MAA & NAB & NAC  |  MAB & NAC  |  MAC  ; 
assign pad = ~PAD;  //complement 
assign KDD = ~kdd;  //complement 
assign KDH = ~kdh;  //complement 
assign HDD =  DDD & cdd  ; 
assign hdd = ~HDD;  //complement  
assign HDE =  DDA & DDB & DDC & DDD  ; 
assign hde = ~HDE;  //complement 
assign KHD = ~khd;  //complement 
assign KHH = ~khh;  //complement 
assign HHD =  DHD & chd  ; 
assign hhd = ~HHD;  //complement  
assign KHC = ~khc;  //complement 
assign KHG = ~khg;  //complement 
assign HHA =  DHA & cha  ; 
assign hha = ~HHA;  //complement 
assign HHB =  DHB & chb  ; 
assign hhb = ~HHB;  //complement 
assign HHC =  DHC & chc  ; 
assign hhc = ~HHC;  //complement 
assign PAH =  QAF & NAE & NAF & NAG  |  MAE & NAF & NAG  |  MAF & NAG  |  MAG  ; 
assign pah = ~PAH;  //complement 
assign ghh =  dha & chb & chc  |  dhb & chc  |  dhc  ; 
assign GHH = ~ghh;  //complement 
assign chc = ~CHC;  //complement 
assign dhc = ~DHC;  //complement 
assign ghf =  dha  ; 
assign GHF = ~ghf;  //complement 
assign ghg =  dha & chb  |  dhb  ; 
assign GHG = ~ghg;  //complement 
assign chd = ~CHD;  //complement 
assign dhd = ~DHD;  //complement 
assign bdc = ~BDC;  //complement 
assign omc = ~OMC;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign QHG = QEG; 
assign qhg = ~QHG; //complement 
assign QHH = QEH; 
assign qhh = ~QHH;  //complement 
assign QIG = QEG; 
assign qig = ~QIG;  //complement 
assign QIH = QEH; 
assign qih = ~QIH;  //complement 
assign bdd = ~BDD;  //complement 
assign omd = ~OMD;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign eah = ~EAH;  //complement 
assign ebh = ~EBH;  //complement 
assign ech = ~ECH;  //complement 
assign edh = ~EDH;  //complement 
assign rao = ~RAO;  //complement 
assign rap = ~RAP;  //complement 
assign aeo = ~AEO;  //complement 
assign aep = ~AEP;  //complement 
assign jic =  sai & saj & sak & sal & sam & san  ; 
assign JIC = ~jic;  //complement  
assign jid =  sam & san & sao & sap  ; 
assign JID = ~jid;  //complement 
assign REO = RAO; 
assign reo = ~REO; //complement 
assign REP = RAP; 
assign rep = ~REP;  //complement 
assign RIO = RAO; 
assign rio = ~RIO;  //complement 
assign RIP = RAP; 
assign rip = ~RIP;  //complement 
assign tld = ~TLD;  //complement 
assign tll = ~TLL;  //complement 
assign tmd = ~TMD;  //complement 
assign tml = ~TML;  //complement 
assign ago = ~AGO;  //complement 
assign agp = ~AGP;  //complement 
assign eeh = ~EEH;  //complement 
assign efh = ~EFH;  //complement 
assign egh = ~EGH;  //complement 
assign ehh = ~EHH;  //complement 
assign RFO = RBO; 
assign rfo = ~RFO; //complement 
assign RFP = RBP; 
assign rfp = ~RFP;  //complement 
assign RJO = RBO; 
assign rjo = ~RJO;  //complement 
assign RJP = RBP; 
assign rjp = ~RJP;  //complement 
assign tlh = ~TLH;  //complement 
assign tlp = ~TLP;  //complement 
assign tmh = ~TMH;  //complement 
assign tmp = ~TMP;  //complement 
assign aio = ~AIO;  //complement 
assign aip = ~AIP;  //complement 
assign EIH = ~eih;  //complement 
assign EJH = ~ejh;  //complement 
assign EKH = ~ekh;  //complement 
assign rbo = ~RBO;  //complement 
assign rbp = ~RBP;  //complement 
assign ako = ~AKO;  //complement 
assign akp = ~AKP;  //complement 
assign ELH = ~elh;  //complement 
assign EPH = ~eph;  //complement 
assign bhc = ~BHC;  //complement 
assign oma = ~OMA;  //complement 
assign amo = ~AMO;  //complement 
assign amp = ~AMP;  //complement 
assign EMH = ~emh;  //complement 
assign ENH = ~enh;  //complement 
assign EOH = ~eoh;  //complement 
assign bhd = ~BHD;  //complement 
assign omb = ~OMB;  //complement 
assign aoo = ~AOO;  //complement 
assign aop = ~AOP;  //complement 
assign jig =  sbi & sbj & sbk & sbl & sbm & sbn  ; 
assign JIG = ~jig;  //complement  
assign jih =  sbm & sbn & sbo & sbp  ; 
assign JIH = ~jih;  //complement 
assign JAO =  AAO & EAH  |  ABO & EBH  |  ACO & ECH  |  ADO & EDH  ; 
assign jao = ~JAO;  //complement 
assign JEO =  AAO & EAH  |  ABO & EBH  |  ACO & ECH  |  ADO & EDH  ; 
assign jeo = ~JEO; //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign rco = ~RCO;  //complement 
assign rgo = ~RGO;  //complement 
assign QEG = ~qeg;  //complement 
assign QEH = ~qeh;  //complement 
assign JAP =  AAP & EAH  |  ABP & EBH  |  ACP & ECH  |  ADP & EDH  ; 
assign jap = ~JAP;  //complement 
assign JEP =  AAP & EAH  |  ABP & EBH  |  ACP & ECH  |  ADP & EDH  ; 
assign jep = ~JEP; //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign rcp = ~RCP;  //complement 
assign rgp = ~RGP;  //complement 
assign oka = ~OKA;  //complement 
assign JBO =  AEO & EEH  |  AFO & EFH  |  AGO & EGH  |  AHO & EHH  ; 
assign jbo = ~JBO;  //complement 
assign JFO =  AEO & EEH  |  AFO & EFH  |  AGO & EGH  |  AHO & EHH  ; 
assign jfo = ~JFO; //complement 
assign afo = ~AFO;  //complement 
assign afp = ~AFP;  //complement 
assign ogo = ~OGO;  //complement 
assign sao = ~SAO;  //complement 
assign sco = ~SCO;  //complement 
assign oao = ~OAO;  //complement 
assign oco = ~OCO;  //complement 
assign oeo = ~OEO;  //complement 
assign JBP =  AEP & EEH  |  AFP & EFH  |  AGP & EGH  |  AHP & EHH  ; 
assign jbp = ~JBP;  //complement 
assign JFP =  AEP & EEH  |  AFP & EFH  |  AGP & EGH  |  AHP & EHH  ; 
assign jfp = ~JFP; //complement 
assign aho = ~AHO;  //complement 
assign ahp = ~AHP;  //complement 
assign ogp = ~OGP;  //complement 
assign sap = ~SAP;  //complement 
assign scp = ~SCP;  //complement 
assign oap = ~OAP;  //complement 
assign ocp = ~OCP;  //complement 
assign oep = ~OEP;  //complement 
assign JCO =  AIO & EIH  |  AJO & EJH  |  AKO & EKH  |  ALO & ELH  ; 
assign jco = ~JCO;  //complement 
assign JGO =  AIO & EIH  |  AJO & EJH  |  AKO & EKH  |  ALO & ELH  ; 
assign jgo = ~JGO; //complement 
assign ajo = ~AJO;  //complement 
assign ajp = ~AJP;  //complement 
assign oho = ~OHO;  //complement 
assign sbo = ~SBO;  //complement 
assign obo = ~OBO;  //complement 
assign odo = ~ODO;  //complement 
assign ofo = ~OFO;  //complement 
assign JCP =  AIP & EIH  |  AJP & EJH  |  AKP & EKH  |  ALP & ELH  ; 
assign jcp = ~JCP;  //complement 
assign JGP =  AIP & EIH  |  AJP & EJH  |  AKP & EKH  |  ALP & ELH  ; 
assign jgp = ~JGP; //complement 
assign alo = ~ALO;  //complement 
assign alp = ~ALP;  //complement 
assign ohp = ~OHP;  //complement 
assign sbp = ~SBP;  //complement 
assign obp = ~OBP;  //complement 
assign odp = ~ODP;  //complement 
assign ofp = ~OFP;  //complement 
assign JDO =  AMO & EMH  |  ANO & ENH  |  AOO & EOH  |  APO & EPH  ; 
assign jdo = ~JDO;  //complement 
assign JHO =  AMO & EMH  |  ANO & ENH  |  AOO & EOH  |  APO & EPH  ; 
assign jho = ~JHO; //complement 
assign ano = ~ANO;  //complement 
assign anp = ~ANP;  //complement 
assign rdo = ~RDO;  //complement 
assign rho = ~RHO;  //complement 
assign qka = ~QKA;  //complement 
assign OLA = ~ola;  //complement 
assign JDP =  AMP & EMH  |  ANP & ENH  |  AOP & EOH  |  APP & EPH  ; 
assign jdp = ~JDP;  //complement 
assign JHP =  AMP & EMH  |  ANP & ENH  |  AOP & EOH  |  APP & EPH  ; 
assign jhp = ~JHP; //complement 
assign apo = ~APO;  //complement 
assign app = ~APP;  //complement 
assign rdp = ~RDP;  //complement 
assign rhp = ~RHP;  //complement 
assign oij = ~OIJ;  //complement 
assign okb = ~OKB;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iff = ~IFF; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
assign ihm = ~IHM; //complement 
assign ihn = ~IHN; //complement 
assign iho = ~IHO; //complement 
assign ihp = ~IHP; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign iic = ~IIC; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ila = ~ILA; //complement 
assign ima = ~IMA; //complement 
always@(posedge IZZ )
   begin 
 CAA <=  BAA & JAA  |  BAA & JBA  ; 
 DAA <=  JAA & JAA  |  JBA & JBA  |  BAA  ; 
 CAB <=  BAB & JAB  |  BAB & JBB  ; 
 DAB <=  JAB & JAB  |  JBB & JBB  |  BAB  ; 
 kaa <=  haa  |  tbe  ; 
 kae <=  HAA  |  tbe  ; 
 kab <=  gab & hab  |  GAB & HAB  |  tbf  ; 
 kaf <=  gaf & hab  |  GAF & HAB  |  tbf  ; 
 maa <= gae ; 
 naa <= hae ; 
 keb <=  geb & heb  |  GEB & HEB  |  tbh  ; 
 kef <=  gef & heb  |  GEF & HEB  |  tbh  ; 
 mae <= gee ; 
 nae <= hee ; 
 kea <=  hea  |  tbg  ; 
 kee <=  HEA  |  tbg  ; 
 CEA <=  BEA & JCA  |  BEA & JDA  ; 
 DEA <=  JCA & JCA  |  JDA & JDA  |  BEA  ; 
 CEB <=  BEB & JCB  |  BEB & JDB  ; 
 DEB <=  JCB & JCB  |  JDB & JDB  |  BEB  ; 
 BAA <=  jaa & jba & tja  |  JAA & TJA  |  JBA & TJC  ; 
 AAA <=  REA & TKA  |  RCA & TKA  |  AAA & tka  ; 
 AAB <=  REB & TKA  |  RCB & TKA  |  AAB & tka  ; 
 BAB <=  jab & jbb & tjb  |  JAB & TJB  |  JBB & TJD  ; 
 ACA <=  REA & TKC  |  RCA & TKC  |  ACA & tkc  ; 
 ACB <=  REB & TKC  |  RCB & TKC  |  ACB & tkc  ; 
 EAA <= qja & QHA ; 
 EBA <= qja & QHB ; 
 ECA <= qja & QHC ; 
 EDA <= qja & QHD ; 
 RAA <=  KAA & paa  |  KAE & PAA  |  LAA & QCB  ; 
 RAB <=  KAB & paa  |  KAF & PAA  |  LAB & QCB  ; 
 AEA <=  REA & TKE  |  RCA & TKE  |  AEA & tke  ; 
 AEB <=  REB & TKE  |  RCB & TKE  |  AEB & tke  ; 
 TAD <= FAD ; 
 TAL <= FAD ; 
 TKD <= FAD ; 
 TKL <= FAD ; 
 AGA <=  REA & TKG  |  RCA & TKG  |  AGA & tkg  ; 
 AGB <=  REB & TKG  |  RCB & TKG  |  AGB & tkg  ; 
 EEA <= qjc & QHE ; 
 EFA <= qjc & QHF ; 
 EGA <= qjc & QHG ; 
 EHA <= qjc & QHH ; 
 TAH <= FAH ; 
 TAP <= FAH ; 
 TKH <= FAH ; 
 TKP <= FAH ; 
 AIA <=  RFA & TAI  |  RDA & TAI  |  AIA & tai  ; 
 AIB <=  RFB & TAI  |  RDB & TAI  |  AIB & tai  ; 
 eia <= ZZI & QJA |  qha & qja ; 
 eja <= ZZI & QJA |  qhb & qja ; 
 eka <= ZZI & QJA |  qhc & qja ; 
 RBA <=  KEA & pae  |  KEE & PAE  ; 
 RBB <=  KEB & pae  |  KEF & PAE  ; 
 AKA <=  RFA & TAK  |  RDA & TAK  |  AKA & tak  ; 
 AKB <=  RFB & TAK  |  RDB & TAK  |  AKB & tak  ; 
 ela <= ZZI & QJI |  qhd & qji ; 
 epa <= ZZI & QJI |  qhh & qji ; 
 BEA <=  jca & jda & tje  |  JCA & TJE  |  JDA & TJG  ; 
 AMA <=  RFA & TAM  |  RDA & TAM  |  AMA & tam  ; 
 AMB <=  RFB & TAM  |  RDB & TAM  |  AMB & tam  ; 
 ema <= ZZI & QJC |  qhe & qjc ; 
 ena <= ZZI & QJC |  qhf & qjc ; 
 eoa <= ZZI & QJC |  qhg & qjc ; 
 BEB <=  jcb & jdb & tjf  |  JCB & TJF  |  JDB & TJH  ; 
 AOA <=  RFA & TAO  |  RDA & TAO  |  AOA & tao  ; 
 AOB <=  RFB & TAO  |  RDB & TAO  |  AOB & tao  ; 
 ABA <=  RIA & TKB  |  RGA & TKB  |  ABA & tkb  ; 
 ABB <=  RIB & TKB  |  RGB & TKB  |  ABB & tkb  ; 
 RCA <=  IAA & TCE  |  ICA & TDE  |  IEA & TEE  |  IGA & TFE  ; 
 RGA <=  IAA & TCE  |  ICA & TDE  |  IEA & TEE  |  IGA & TFE  ; 
 laa <=  jea & jfa & QFB  |  laa & qfb  ; 
 oja <=  jea & jfa & QFB  |  laa & qfb  ; 
 ADA <=  RIA & TKD  |  RGA & TKD  |  ADA & tkd  ; 
 ADB <=  RIB & TKD  |  RGB & TKD  |  ADB & tkd  ; 
 RCB <=  IAB & TCF  |  ICB & TDF  |  IEB & TEF  |  IGB & TFF  ; 
 RGB <=  IAB & TCF  |  ICB & TDF  |  IEB & TEF  |  IGB & TFF  ; 
 lab <=  jeb & jfb & QFC  |  lab & qfc  ; 
 ojb <=  jeb & jfb & QFC  |  lab & qfc  ; 
 AFA <=  RIA & TKF  |  RGA & TKF  |  AFA & tkf  ; 
 AFB <=  RIB & TKF  |  RGB & TKF  |  AFB & tkf  ; 
 OGA <=  JEA  |  JFA  ; 
 OIA <=  JEA  |  JFA  ; 
 SAA <=  JEA  |  JFA  ; 
 OAA <=  JEA  |  JFA  ; 
 OCA <=  JEA  |  JFA  ; 
 OEA <=  JEA  |  JFA  ; 
 AHA <=  RIA & TKH  |  RGA & TKH  |  AHA & tkh  ; 
 AHB <=  RIB & TKH  |  RGB & TKH  |  AHB & tkh  ; 
 OGB <=  JEB  |  JFB  ; 
 OIB <=  JEB  |  JFB  ; 
 SAB <=  JEB  |  JFB  ; 
 OAB <=  JEB  |  JFB  ; 
 OCB <=  JEB  |  JFB  ; 
 OEB <=  JEB  |  JFB  ; 
 AJA <=  RJA & TAJ  |  RHA & TAJ  |  AJA & taj  ; 
 AJB <=  RJB & TAJ  |  RHB & TAJ  |  AJB & taj  ; 
 OHA <=  JGA  |  JHA  ; 
 SBA <=  JGA  |  JHA  ; 
 OBA <=  JGA  |  JHA  ; 
 ODA <=  JGA  |  JHA  ; 
 OFA <=  JGA  |  JHA  ; 
 ALA <=  RJA & TAL  |  RHA & TAL  |  ALA & tal  ; 
 ALB <=  RJB & TAL  |  RHB & TAL  |  ALB & tal  ; 
 OHB <=  JGB  |  JHB  ; 
 SBB <=  JGB  |  JHB  ; 
 OBB <=  JGB  |  JHB  ; 
 ODB <=  JGB  |  JHB  ; 
 OFB <=  JGB  |  JHB  ; 
 ANA <=  RJA & TAN  |  RHA & TAN  |  ANA & tan  ; 
 ANB <=  RJB & TAN  |  RHB & TAN  |  ANB & tan  ; 
 RDA <=  IBA & TCG  |  IDA & TDG  |  IFA & TEG  |  IHA & TFG  ; 
 RHA <=  IBA & TCG  |  IDA & TDG  |  IFA & TEG  |  IHA & TFG  ; 
 CIA <=  QKA & QFH  |  QAA & QFH  ; 
 APA <=  RJA & TAP  |  RHA & TAP  |  APA & tap  ; 
 APB <=  RJB & TAP  |  RHB & TAP  |  APB & tap  ; 
 RDB <=  IBB & TCH  |  IDB & TDH  |  IFB & TEH  |  IHB & TFH  ; 
 RHB <=  IBB & TCH  |  IDB & TDH  |  IFB & TEH  |  IHB & TFH  ; 
 CAC <=  BAC & JAC  |  BAC & JBC  ; 
 DAC <=  JAC & JAC  |  JBC & JBC  |  BAC  ; 
 CAD <=  BAD & JAD  |  BAD & JBD  ; 
 DAD <=  JAD & JAD  |  JBD & JBD  |  BAD  ; 
 kac <=  gac & hac  |  GAC & HAC  |  tbe  ; 
 kag <=  gag & hac  |  GAG & HAC  |  tbe  ; 
 kad <=  gad & had  |  GAD & HAD  |  tbf  ; 
 kah <=  gah & had  |  GAH & HAD  |  tbf  ; 
 ked <=  ged & hed  |  GED & HED  |  tbh  ; 
 keh <=  geh & hed  |  GEH & HED  |  tbh  ; 
 TAG <= FAG ; 
 TAO <= FAG ; 
 TKG <= FAG ; 
 TKO <= FAG ; 
 kec <=  gec & hec  |  GEC & HEC  |  tbg  ; 
 keg <=  geg & hec  |  GEG & HEC  |  tbg  ; 
 CEC <=  BEC & JCC  |  BEC & JDC  ; 
 DEC <=  JCC & JCC  |  JDC & JDC  |  BEC  ; 
 CED <=  BED & JCD  |  BED & JDD  ; 
 DED <=  JCD & JCD  |  JDD & JDD  |  BED  ; 
 BAC <=  jac & jbc & tja  |  JAC & TJA  |  JBC & TJC  ; 
 AAC <=  REC & TKA  |  RCC & TKA  |  AAC & tka  ; 
 AAD <=  RED & TKA  |  RCD & TKA  |  AAD & tka  ; 
 BAD <=  jad & jbd & tjb  |  JAD & TJB  |  JBD & TJD  ; 
 ACC <=  REC & TKC  |  RCC & TKC  |  ACC & tkc  ; 
 ACD <=  RED & TKC  |  RCD & TKC  |  ACD & tkc  ; 
 EAB <= qjb & QHA ; 
 EBB <= qjb & QHB ; 
 ECB <= qjb & QHC ; 
 EDB <= qjb & QHD ; 
 RAC <=  KAC & paa  |  KAG & PAA  |  LAC & QCB  ; 
 RAD <=  KAD & paa  |  KAH & PAA  |  LAD & QCB  ; 
 AEC <=  REC & TKE  |  RCC & TKE  |  AEC & tke  ; 
 AED <=  RED & TKE  |  RCD & TKE  |  AED & tke  ; 
 TAC <= FAC ; 
 TAK <= FAC ; 
 TKC <= FAC ; 
 TKK <= FAC ; 
 AGC <=  REC & TKG  |  RCC & TKG  |  AGC & tkg  ; 
 AGD <=  RED & TKG  |  RCD & TKG  |  AGD & tkg  ; 
 EEB <= qjd & QHE ; 
 EFB <= qjd & QHF ; 
 EGB <= qjd & QHG ; 
 EHB <= qjd & QHH ; 
 AIC <=  RFC & TAI  |  RDC & TAI  |  AIC & tai  ; 
 AID <=  RFD & TAI  |  RDD & TAI  |  AID & tai  ; 
 eib <= ZZI & QJB |  qha & qjb ; 
 ejb <= ZZI & QJB |  qhb & qjb ; 
 ekb <= ZZI & QJB |  qhc & qjb ; 
 RBC <=  KEC & pae  |  KEG & PAE  ; 
 RBD <=  KED & pae  |  KEH & PAE  ; 
 AKC <=  RFC & TAK  |  RDC & TAK  |  AKC & tak  ; 
 AKD <=  RFD & TAK  |  RDD & TAK  |  AKD & tak  ; 
 elb <= ZZI & QJJ |  qhd & qjj ; 
 epb <= ZZI & QJJ |  qhh & qjj ; 
 BEC <=  jcc & jdc & tje  |  JCC & TJE  |  JDC & TJG  ; 
 AMC <=  RFC & TAM  |  RDC & TAM  |  AMC & tam  ; 
 AMD <=  RFD & TAM  |  RDD & TAM  |  AMD & tam  ; 
 emb <= ZZI & QJD |  qhe & qjd ; 
 enb <= ZZI & QJD |  qhf & qjd ; 
 eob <= ZZI & QJD |  qhg & qjd ; 
 BED <=  jcd & jdd & tjf  |  JCD & TJF  |  JDD & TJH  ; 
 AOC <=  RFC & TAO  |  RDC & TAO  |  AOC & tao  ; 
 AOD <=  RFD & TAO  |  RDD & TAO  |  AOD & tao  ; 
 ABC <=  RIC & TKB  |  RGC & TKB  |  ABC & tkb  ; 
 ABD <=  RID & TKB  |  RGD & TKB  |  ABD & tkb  ; 
 RCC <=  IAC & TCE  |  ICC & TDE  |  IEC & TEE  |  IGC & TFE  ; 
 RGC <=  IAC & TCE  |  ICC & TDE  |  IEC & TEE  |  IGC & TFE  ; 
 lac <=  jec & jfc & QFB  |  lac & qfb  ; 
 ojc <=  jec & jfc & QFB  |  lac & qfb  ; 
 ADC <=  RIC & TKD  |  RGC & TKD  |  ADC & tkd  ; 
 ADD <=  RID & TKD  |  RGD & TKD  |  ADD & tkd  ; 
 RCD <=  IAD & TCF  |  ICD & TDF  |  IED & TEF  |  IGD & TFF  ; 
 RGD <=  IAD & TCF  |  ICD & TDF  |  IED & TEF  |  IGD & TFF  ; 
 lad <=  jed & jfd & QFC  |  lad & qfc  ; 
 ojd <=  jed & jfd & QFC  |  lad & qfc  ; 
 AFC <=  RIC & TKF  |  RGC & TKF  |  AFC & tkf  ; 
 AFD <=  RID & TKF  |  RGD & TKF  |  AFD & tkf  ; 
 OGC <=  JEC  |  JFC  ; 
 OIC <=  JEC  |  JFC  ; 
 SAC <=  JEC  |  JFC  ; 
 OAC <=  JEC  |  JFC  ; 
 OCC <=  JEC  |  JFC  ; 
 OEC <=  JEC  |  JFC  ; 
 AHC <=  RIC & TKH  |  RGC & TKH  |  AHC & tkh  ; 
 AHD <=  RID & TKH  |  RGD & TKH  |  AHD & tkh  ; 
 OGD <=  JED  |  JFD  ; 
 OID <=  JED  |  JFD  ; 
 SAD <=  JED  |  JFD  ; 
 OAD <=  JED  |  JFD  ; 
 OCD <=  JED  |  JFD  ; 
 OED <=  JED  |  JFD  ; 
 AJC <=  RJC & TAJ  |  RHC & TAJ  |  AJC & taj  ; 
 AJD <=  RJD & TAJ  |  RHD & TAJ  |  AJD & taj  ; 
 OHC <=  JGC  |  JHC  ; 
 SBC <=  JGC  |  JHC  ; 
 OBC <=  JGC  |  JHC  ; 
 ODC <=  JGC  |  JHC  ; 
 OFC <=  JGC  |  JHC  ; 
 ALC <=  RJC & TAL  |  RHC & TAL  |  ALC & tal  ; 
 ALD <=  RJD & TAL  |  RHD & TAL  |  ALD & tal  ; 
 OHD <=  JGD  |  JHD  ; 
 SBD <=  JGD  |  JHD  ; 
 OBD <=  JGD  |  JHD  ; 
 ODD <=  JGD  |  JHD  ; 
 OFD <=  JGD  |  JHD  ; 
 ANC <=  RJC & TAN  |  RHC & TAN  |  ANC & tan  ; 
 AND <=  RJD & TAN  |  RHD & TAN  |  AND & tan  ; 
 RDC <=  IBC & TCG  |  IDC & TDG  |  IFC & TEG  |  IHC & TFG  ; 
 RHC <=  IBC & TCG  |  IDC & TDG  |  IFC & TEG  |  IHC & TFG  ; 
 OME <=  RJP & TLB  |  RHP & TLB  |  AJP & tlb  ; 
 APC <=  RJC & TAP  |  RHC & TAP  |  APC & tap  ; 
 APD <=  RJD & TAP  |  RHD & TAP  |  APD & tap  ; 
 RDD <=  IBD & TCH  |  IDD & TDH  |  IFD & TEH  |  IHD & TFH  ; 
 RHD <=  IBD & TCH  |  IDD & TDH  |  IFD & TEH  |  IHD & TFH  ; 
 OMF <=  RJP & TLD  |  RHP & TLD  |  ALP & tld  ; 
 CBA <=  BBA & JAE  |  BBA & JBE  ; 
 DBA <=  JAE & JAE  |  JBE & JBE  |  BBA  ; 
 CBB <=  BBB & JAF  |  BBB & JBF  ; 
 DBB <=  JAF & JAF  |  JBF & JBF  |  BBB  ; 
 kba <=  hba  |  tbe  ; 
 kbe <=  HBA  |  tbe  ; 
 kbb <=  gbb & hbb  |  GBB & HBB  |  tbf  ; 
 kbf <=  gbf & hbb  |  GBF & HBB  |  tbf  ; 
 mab <= gbe ; 
 nab <= hbe ; 
 kfb <=  gfb & hfb  |  GFB & HFB  |  tbh  ; 
 kff <=  gff & hfb  |  GFF & HFB  |  tbh  ; 
 maf <= gfe ; 
 naf <= hfe ; 
 kfa <=  hfa  |  tbg  ; 
 kfe <=  HFA  |  tbg  ; 
 OMG <=  RJP & TLF  |  RHP & TLF  |  ANP & tlf  ; 
 CFA <=  BFA & JCE  |  BFA & JDE  ; 
 DFA <=  JCE & JCE  |  JDE & JDE  |  BFA  ; 
 OMH <=  RJP & TLH  |  RHP & TLH  |  APP & tlh  ; 
 CFB <=  BFB & JCF  |  BFB & JDF  ; 
 DFB <=  JCF & JCF  |  JDF & JDF  |  BFB  ; 
 BBA <=  jae & jbe & tja  |  JAE & TJA  |  JBE & TJC  ; 
 AAE <=  REE & TKI  |  RCE & TKI  |  AAE & tki  ; 
 AAF <=  REF & TKI  |  RCF & TKI  |  AAF & tki  ; 
 BBB <=  jaf & jbf & tjb  |  JAF & TJB  |  JBF & TJD  ; 
 ACE <=  REE & TKK  |  RCE & TKK  |  ACE & tkk  ; 
 ACF <=  REF & TKK  |  RCF & TKK  |  ACF & tkk  ; 
 EAC <= qja & QHA ; 
 EBC <= qja & QHB ; 
 ECC <= qja & QHC ; 
 EDC <= qja & QHD ; 
 RAE <=  KBA & pab  |  KBE & PAB  |  LAE & QCB  ; 
 RAF <=  KBB & pab  |  KBF & PAB  |  LAF & QCB  ; 
 AEE <=  REE & TKM  |  RCE & TKM  |  AEE & tkm  ; 
 AEF <=  REF & TKM  |  RCF & TKM  |  AEF & tkm  ; 
 TAB <= FAB ; 
 TAJ <= FAB ; 
 TKB <= FAB ; 
 TKJ <= FAB ; 
 AGE <=  REE & TKO  |  RCE & TKO  |  AGE & tko  ; 
 AGF <=  REF & TKO  |  RCF & TKO  |  AGF & tko  ; 
 EEC <= qjc & QHE ; 
 EFC <= qjc & QHF ; 
 EGC <= qjc & QHG ; 
 EHC <= qjc & QHH ; 
 TAF <= FAF ; 
 TAN <= FAF ; 
 TKF <= FAF ; 
 TKN <= FAF ; 
 AIE <=  RFE & TAA  |  RDE & TAA  |  AIE & taa  ; 
 AIF <=  RFF & TAA  |  RDF & TAA  |  AIF & taa  ; 
 eic <= ZZI & QJA |  qha & qja ; 
 ejc <= ZZI & QJA |  qhb & qja ; 
 ekc <= ZZI & QJA |  qhc & qja ; 
 RBE <=  KFA & paf  |  KFE & PAF  ; 
 RBF <=  KFB & paf  |  KFF & PAF  ; 
 AKE <=  RFE & TAC  |  RDE & TAC  |  AKE & tac  ; 
 AKF <=  RFF & TAC  |  RDF & TAC  |  AKF & tac  ; 
 elc <= ZZI & QJI |  qhd & qji ; 
 epc <= ZZI & QJI |  qhh & qji ; 
 BFA <=  jce & jde & tje  |  JCE & TJE  |  JDE & TJG  ; 
 AME <=  RFE & TAE  |  RDE & TAE  |  AME & tae  ; 
 AMF <=  RFF & TAE  |  RDF & TAE  |  AMF & tae  ; 
 emc <= ZZI & QJC |  qhe & qjc ; 
 enc <= ZZI & QJC |  qhf & qjc ; 
 eoc <= ZZI & QJC |  qhg & qjc ; 
 BFB <=  jcf & jdf & tjf  |  JCF & TJF  |  JDF & TJH  ; 
 AOE <=  RFE & TAG  |  RDE & TAG  |  AOE & tag  ; 
 AOF <=  RFF & TAG  |  RDF & TAG  |  AOF & tag  ; 
 ABE <=  RIE & TKJ  |  RGE & TKJ  |  ABE & tkj  ; 
 ABF <=  RIF & TKJ  |  RGF & TKJ  |  ABF & tkj  ; 
 RCE <=  IAE & TCE  |  ICE & TDE  |  IEE & TEE  |  IGE & TFE  ; 
 RGE <=  IAE & TCE  |  ICE & TDE  |  IEE & TEE  |  IGE & TFE  ; 
 lae <=  jee & jfe & QFB  |  lae & qfb  ; 
 oje <=  jee & jfe & QFB  |  lae & qfb  ; 
 ADE <=  RIE & TKL  |  RGE & TKL  |  ADE & tkl  ; 
 ADF <=  RIF & TKL  |  RGF & TKL  |  ADF & tkl  ; 
 RCF <=  IAF & TCF  |  ICF & TDF  |  IEF & TEF  |  IGF & TFF  ; 
 RGF <=  IAF & TCF  |  ICF & TDF  |  IEF & TEF  |  IGF & TFF  ; 
 laf <=  jef & jff & QFC  |  laf & qfc  ; 
 ojf <=  jef & jff & QFC  |  laf & qfc  ; 
 AFE <=  RIE & TKN  |  RGE & TKN  |  AFE & tkn  ; 
 AFF <=  RIF & TKN  |  RGF & TKN  |  AFF & tkn  ; 
 OGE <=  JEE  |  JFE  ; 
 OIE <=  JEE  |  JFE  ; 
 SAE <=  JEE  |  JFE  ; 
 OAE <=  JEE  |  JFE  ; 
 OCE <=  JEE  |  JFE  ; 
 OEE <=  JEE  |  JFE  ; 
 AHE <=  RIE & TKP  |  RGE & TKP  |  AHE & tkp  ; 
 AHF <=  RIF & TKP  |  RGF & TKP  |  AHF & tkp  ; 
 OGF <=  JEF  |  JFF  ; 
 OIF <=  JEF  |  JFF  ; 
 SAF <=  JEF  |  JFF  ; 
 OAF <=  JEF  |  JFF  ; 
 OCF <=  JEF  |  JFF  ; 
 OEF <=  JEF  |  JFF  ; 
 AJE <=  RJE & TAB  |  RHE & TAB  |  AJE & tab  ; 
 AJF <=  RJF & TAB  |  RHF & TAB  |  AJF & tab  ; 
 OHE <=  JGE  |  JHE  ; 
 SBE <=  JGE  |  JHE  ; 
 OBE <=  JGE  |  JHE  ; 
 ODE <=  JGE  |  JHE  ; 
 OFE <=  JGE  |  JHE  ; 
 ALE <=  RJE & TAD  |  RHE & TAD  |  ALE & tad  ; 
 ALF <=  RJF & TAD  |  RHF & TAD  |  ALF & tad  ; 
 OHF <=  JGF  |  JHF  ; 
 SBF <=  JGF  |  JHF  ; 
 OBF <=  JGF  |  JHF  ; 
 ODF <=  JGF  |  JHF  ; 
 OFF <=  JGF  |  JHF  ; 
 ANE <=  RJE & TAF  |  RHE & TAF  |  ANE & taf  ; 
 ANF <=  RJF & TAF  |  RHF & TAF  |  ANF & taf  ; 
 RDE <=  IBE & TCG  |  IDE & TDG  |  IFE & TEG  |  IHE & TFG  ; 
 RHE <=  IBE & TCG  |  IDE & TDG  |  IFE & TEG  |  IHE & TFG  ; 
 APE <=  RJE & TAH  |  RHE & TAH  |  APE & tah  ; 
 APF <=  RJF & TAH  |  RHF & TAH  |  APF & tah  ; 
 RDF <=  IBF & TCH  |  IDF & TDH  |  IFF & TEH  |  IHF & TFH  ; 
 RHF <=  IBF & TCH  |  IDF & TDH  |  IFF & TEH  |  IHF & TFH  ; 
 CBC <=  BBC & JAG  |  BBC & JBG  ; 
 DBC <=  JAG & JAG  |  JBG & JBG  |  BBC  ; 
 CBD <=  BBD & JAH  |  BBD & JBH  ; 
 DBD <=  JAH & JAH  |  JBH & JBH  |  BBD  ; 
 kbc <=  gbc & hbc  |  GBC & HBC  |  tbe  ; 
 kbg <=  gbg & hbc  |  GBG & HBC  |  tbe  ; 
 kbd <=  gbd & hbd  |  GBD & HBD  |  tbf  ; 
 kbh <=  gbh & hbd  |  GBH & HBD  |  tbf  ; 
 TJA <= qaa ; 
 TJB <= qaa ; 
 TJC <= qaa ; 
 TJD <= qaa ; 
 kfd <=  gfd & hfd  |  GFD & HFD  |  tbh  ; 
 kfh <=  gfh & hfd  |  GFH & HFD  |  tbh  ; 
 TJE <= qaa ; 
 TJF <= qaa ; 
 TJG <= qaa ; 
 TJH <= qaa ; 
 kfc <=  gfc & hfc  |  GFC & HFC  |  tbg  ; 
 kfg <=  gfg & hfc  |  GFG & HFC  |  tbg  ; 
 CFC <=  BFC & JCG  |  BFC & JDG  ; 
 DFC <=  JCG & JCG  |  JDG & JDG  |  BFC  ; 
 CFD <=  BFD & JCH  |  BFD & JDH  ; 
 DFD <=  JCH & JCH  |  JDH & JDH  |  BFD  ; 
 BBC <=  jag & jbg & tja  |  JAG & TJA  |  JBG & TJC  ; 
 AAG <=  REG & TKI  |  RCG & TKI  |  AAG & tki  ; 
 AAH <=  REH & TKI  |  RCH & TKI  |  AAH & tki  ; 
 qfe <=  ikb  |  ila  ; 
 qff <=  ikb  |  ila  ; 
 qfg <=  ikb  |  ila  ; 
 BBD <=  jah & jbh & tjb  |  JAH & TJB  |  JBH & TJD  ; 
 ACG <=  REG & TKK  |  RCG & TKK  |  ACG & tkk  ; 
 ACH <=  REH & TKK  |  RCH & TKK  |  ACH & tkk  ; 
 EAD <= qjb & QHA ; 
 EBD <= qjb & QHB ; 
 ECD <= qjb & QHC ; 
 EDD <= qjb & QHD ; 
 RAG <=  KBC & pab  |  KBG & PAB  ; 
 RAH <=  KBD & pab  |  KBH & PAB  ; 
 AEG <=  REG & TKM  |  RCG & TKM  |  AEG & tkm  ; 
 AEH <=  REH & TKM  |  RCH & TKM  |  AEH & tkm  ; 
 QFB <= qbb & QFA ; 
 QFC <= qbb & QFA ; 
 TAA <= FAA ; 
 TAI <= FAA ; 
 TKA <= FAA ; 
 TKI <= FAA ; 
 AGG <=  REG & TKO  |  RCG & TKO  |  AGG & tko  ; 
 AGH <=  REH & TKO  |  RCH & TKO  |  AGH & tko  ; 
 EED <= qjd & QHE ; 
 EFD <= qjd & QHF ; 
 EGD <= qjd & QHG ; 
 EHD <= qjd & QHH ; 
 TAE <= FAE ; 
 TAM <= FAE ; 
 TKE <= FAE ; 
 TKM <= FAE ; 
 AIG <=  RFG & TAA  |  RDG & TAA  |  AIG & taa  ; 
 AIH <=  RFH & TAA  |  RDH & TAA  |  AIH & taa  ; 
 eid <= ZZI & QJB |  qha & qjb ; 
 ejd <= ZZI & QJB |  qhb & qjb ; 
 ekd <= ZZI & QJB |  qhc & qjb ; 
 RBG <=  KFC & paf  |  KFG & PAF  ; 
 RBH <=  KFD & paf  |  KFH & PAF  ; 
 AKG <=  RFG & TAC  |  RDG & TAC  |  AKG & tac  ; 
 AKH <=  RFH & TAC  |  RDH & TAC  |  AKH & tac  ; 
 eld <= ZZI & QJJ |  qhd & qjj ; 
 epd <= ZZI & QJJ |  qhh & qjj ; 
 BFC <=  jcg & jdg & tje  |  JCG & TJE  |  JDG & TJG  ; 
 AMG <=  RFG & TAE  |  RDG & TAE  |  AMG & tae  ; 
 AMH <=  RFH & TAE  |  RDH & TAE  |  AMH & tae  ; 
 emd <= ZZI & QJD |  qhe & qjd ; 
 end <= ZZI & QJD |  qhf & qjd ; 
 eod <= ZZI & QJD |  qhg & qjd ; 
 BFD <=  jch & jdh & tjf  |  JCH & TJF  |  JDH & TJH  ; 
 AOG <=  RFG & TAG  |  RDG & TAG  |  AOG & tag  ; 
 AOH <=  RFH & TAG  |  RDH & TAG  |  AOH & tag  ; 
 TBE <= QBC ; 
 TBF <= QBC ; 
 TBG <= QBC ; 
 TBH <= QBC ; 
 ABG <=  RIG & TKJ  |  RGG & TKJ  |  ABG & tkj  ; 
 ABH <=  RIH & TKJ  |  RGH & TKJ  |  ABH & tkj  ; 
 RCG <=  IAG & TCE  |  ICG & TDE  |  IEG & TEE  |  IGG & TFE  ; 
 RGG <=  IAG & TCE  |  ICG & TDE  |  IEG & TEE  |  IGG & TFE  ; 
 ADG <=  RIG & TKL  |  RGG & TKL  |  ADG & tkl  ; 
 ADH <=  RIH & TKL  |  RGH & TKL  |  ADH & tkl  ; 
 RCH <=  IAH & TCF  |  ICH & TDF  |  IEH & TEF  |  IGH & TFF  ; 
 RGH <=  IAH & TCF  |  ICH & TDF  |  IEH & TEF  |  IGH & TFF  ; 
 AFG <=  RIG & TKN  |  RGG & TKN  |  AFG & tkn  ; 
 AFH <=  RIH & TKN  |  RGH & TKN  |  AFH & tkn  ; 
 OGG <=  JEG  |  JFG  ; 
 OIG <=  JEG  |  JFG  ; 
 SAG <=  JEG  |  JFG  ; 
 OAG <=  JEG  |  JFG  ; 
 OCG <=  JEG  |  JFG  ; 
 OEG <=  JEG  |  JFG  ; 
 AHG <=  RIG & TKP  |  RGG & TKP  |  AHG & tkp  ; 
 AHH <=  RIH & TKP  |  RGH & TKP  |  AHH & tkp  ; 
 OGH <=  JEH  |  JFH  ; 
 OIH <=  JEH  |  JFH  ; 
 SAH <=  JEH  |  JFH  ; 
 OAH <=  JEH  |  JFH  ; 
 OCH <=  JEH  |  JFH  ; 
 OEH <=  JEH  |  JFH  ; 
 AJG <=  RJG & TAB  |  RHG & TAB  |  AJG & tab  ; 
 AJH <=  RJH & TAB  |  RHH & TAB  |  AJH & tab  ; 
 OHG <=  JGG  |  JHG  ; 
 SBG <=  JGG  |  JHG  ; 
 OBG <=  JGG  |  JHG  ; 
 ODG <=  JGG  |  JHG  ; 
 OFG <=  JGG  |  JHG  ; 
 ALG <=  RJG & TAD  |  RHG & TAD  |  ALG & tad  ; 
 ALH <=  RJH & TAD  |  RHH & TAD  |  ALH & tad  ; 
 OHH <=  JGH  |  JHH  ; 
 SBH <=  JGH  |  JHH  ; 
 OBH <=  JGH  |  JHH  ; 
 ODH <=  JGH  |  JHH  ; 
 OFH <=  JGH  |  JHH  ; 
 ANG <=  RJG & TAF  |  RHG & TAF  |  ANG & taf  ; 
 ANH <=  RJH & TAF  |  RHH & TAF  |  ANH & taf  ; 
 RDG <=  IBG & TCG  |  IDG & TDG  |  IFG & TEG  |  IHG & TFG  ; 
 RHG <=  IBG & TCG  |  IDG & TDG  |  IFG & TEG  |  IHG & TFG  ; 
 APG <=  RJG & TAH  |  RHG & TAH  |  APG & tah  ; 
 APH <=  RJH & TAH  |  RHH & TAH  |  APH & tah  ; 
 RDH <=  IBH & TCH  |  IDH & TDH  |  IFH & TEH  |  IHH & TFH  ; 
 RHH <=  IBH & TCH  |  IDH & TDH  |  IFH & TEH  |  IHH & TFH  ; 
 CCA <=  BCA & JAI  |  BCA & JBI  ; 
 DCA <=  JAI & JAI  |  JBI & JBI  |  BCA  ; 
 CCB <=  BCB & JAJ  |  BCB & JBJ  ; 
 DCB <=  JAJ & JAJ  |  JBJ & JBJ  |  BCB  ; 
 kca <=  hca  |  tba  ; 
 kce <=  HCA  |  tba  ; 
 TIA <= qaa ; 
 TIB <= qaa ; 
 TIC <= qaa ; 
 TID <= qaa ; 
 kcb <=  gcb & hcb  |  GCB & HCB  |  tbb  ; 
 kcf <=  gcf & hcb  |  GCF & HCB  |  tbb  ; 
 mac <= gce ; 
 nac <= hce ; 
 kgb <=  ggb & hgb  |  GGB & HGB  |  tbd  ; 
 kgf <=  ggf & hgb  |  GGF & HGB  |  tbd  ; 
 mag <= gge ; 
 nag <= hge ; 
 kga <=  hga  |  tbc  ; 
 kge <=  HGA  |  tbc  ; 
 TIE <= qaa ; 
 TIF <= qaa ; 
 TIG <= qaa ; 
 TIH <= qaa ; 
 CGA <=  BGA & JCI  |  BGA & JDI  ; 
 DGA <=  JCI & JCI  |  JDI & JDI  |  BGA  ; 
 CGB <=  BGB & JCJ  |  BGB & JDJ  ; 
 DGB <=  JCJ & JCJ  |  JDJ & JDJ  |  BGB  ; 
 BCA <=  jai & jbi & tia  |  JAI & TIA  |  JBI & TIC  ; 
 AAI <=  REI & TMA  |  RCI & TMA  |  AAI & tma  ; 
 AAJ <=  REJ & TMA  |  RCJ & TMA  |  AAJ & tma  ; 
 BCB <=  jaj & jbj & tib  |  JAJ & TIB  |  JBJ & TID  ; 
 ACI <=  REI & TMC  |  RCI & TMC  |  ACI & tmc  ; 
 ACJ <=  REJ & TMC  |  RCJ & TMC  |  ACJ & tmc  ; 
 EAE <= qja & QIA ; 
 EBE <= qja & QIB ; 
 ECE <= qja & QIC ; 
 EDE <= qja & QID ; 
 RAI <=  KCA & pac  |  KCE & PAC  ; 
 RAJ <=  KCB & pac  |  KCF & PAC  ; 
 AEI <=  REI & TME  |  RCI & TME  |  AEI & tme  ; 
 AEJ <=  REJ & TME  |  RCJ & TME  |  AEJ & tme  ; 
 QAB <= QAA ; 
 QAC <= QAB ; 
 QAD <= QAC ; 
 TLA <= FBA ; 
 TLI <= FBA ; 
 TMA <= FBA ; 
 TMI <= FBA ; 
 AGI <=  REI & TMG  |  RCI & TMG  |  AGI & tmg  ; 
 AGJ <=  REJ & TMG  |  RCJ & TMG  |  AGJ & tmg  ; 
 EEE <= qjc & QIE ; 
 EFE <= qjc & QIF ; 
 EGE <= qjc & QIG ; 
 EHE <= qjc & QIH ; 
 TLE <= FBE ; 
 TLM <= FBE ; 
 TME <= FBE ; 
 TMM <= FBE ; 
 AII <=  RFI & TLI  |  RDI & TLI  |  AII & tli  ; 
 AIJ <=  RFJ & TLI  |  RDJ & TLI  |  AIJ & tli  ; 
 eie <= ZZI & QJA |  qia & qja ; 
 eje <= ZZI & QJA |  qib & qja ; 
 eke <= ZZI & QJA |  qic & qja ; 
 RBI <=  KGA & pag  |  KGE & PAG  ; 
 RBJ <=  KGB & pag  |  KGF & PAG  ; 
 AKI <=  RFI & TLK  |  RDI & TLK  |  AKI & tlk  ; 
 AKJ <=  RFJ & TLK  |  RDJ & TLK  |  AKJ & tlk  ; 
 ele <= ZZI & QJI |  qid & qji ; 
 epe <= ZZI & QJI |  qih & qji ; 
 BGA <=  jci & jdi & tie  |  JCI & TIE  |  JDI & TIG  ; 
 AMI <=  RFI & TLM  |  RDI & TLM  |  AMI & tlm  ; 
 AMJ <=  RFJ & TLM  |  RDJ & TLM  |  AMJ & tlm  ; 
 eme <= ZZI & QJC |  qie & qjc ; 
 ene <= ZZI & QJC |  qif & qjc ; 
 eoe <= ZZI & QJC |  qig & qjc ; 
 BGB <=  jcj & jdj & tif  |  JCJ & TIF  |  JDJ & TIH  ; 
 AOI <=  RFI & TLO  |  RDI & TLO  |  AOI & tlo  ; 
 AOJ <=  RFJ & TLO  |  RDJ & TLO  |  AOJ & tlo  ; 
 TBA <= QBC ; 
 TBB <= QBC ; 
 TBC <= QBC ; 
 TBD <= QBC ; 
 ABI <=  RII & TMB  |  RGI & TMB  |  ABI & tmb  ; 
 ABJ <=  RIJ & TMB  |  RGJ & TMB  |  ABJ & tmb  ; 
 RCI <=  IAI & TCA  |  ICI & TDA  |  IEI & TEA  |  IGI & TFA  ; 
 RGI <=  IAI & TCA  |  ICI & TDA  |  IEI & TEA  |  IGI & TFA  ; 
 qea <=  IIC  |  IIB  |  IIA  ; 
 qeb <=  IIC  |  IIB  |  iia  ; 
 ADI <=  RII & TMD  |  RGI & TMD  |  ADI & tmd  ; 
 ADJ <=  RIJ & TMD  |  RGJ & TMD  |  ADJ & tmd  ; 
 RCJ <=  IAJ & TCB  |  ICJ & TDB  |  IEJ & TEB  |  IGJ & TFB  ; 
 RGJ <=  IAJ & TCB  |  ICJ & TDB  |  IEJ & TEB  |  IGJ & TFB  ; 
 QAA <= IKA ; 
 QFA <= ILA ; 
 QFH <= ILA ; 
 AFI <=  RII & TMF  |  RGI & TMF  |  AFI & tmf  ; 
 AFJ <=  RIJ & TMF  |  RGJ & TMF  |  AFJ & tmf  ; 
 OGI <=  JEI  |  JFI  ; 
 SAI <=  JEI  |  JFI  ; 
 OAI <=  JEI  |  JFI  ; 
 OCI <=  JEI  |  JFI  ; 
 OEI <=  JEI  |  JFI  ; 
 AHI <=  RII & TMH  |  RGI & TMH  |  AHI & tmh  ; 
 AHJ <=  RIJ & TMH  |  RGJ & TMH  |  AHJ & tmh  ; 
 OGJ <=  JEJ  |  JFJ  ; 
 SAJ <=  JEJ  |  JFJ  ; 
 OAJ <=  JEJ  |  JFJ  ; 
 OCJ <=  JEJ  |  JFJ  ; 
 OEJ <=  JEJ  |  JFJ  ; 
 AJI <=  RJI & TLJ  |  RHI & TLJ  |  AJI & tlj  ; 
 AJJ <=  RJJ & TLJ  |  RHJ & TLJ  |  AJJ & tlj  ; 
 OHI <=  JGI  |  JHI  ; 
 SBI <=  JGI  |  JHI  ; 
 OBI <=  JGI  |  JHI  ; 
 ODI <=  JGI  |  JHI  ; 
 OFI <=  JGI  |  JHI  ; 
 ALI <=  RJI & TLL  |  RHI & TLL  |  ALI & tll  ; 
 ALJ <=  RJJ & TLL  |  RHJ & TLL  |  ALJ & tll  ; 
 OHJ <=  JGJ  |  JHJ  ; 
 SBJ <=  JGJ  |  JHJ  ; 
 OBJ <=  JGJ  |  JHJ  ; 
 ODJ <=  JGJ  |  JHJ  ; 
 OFJ <=  JGJ  |  JHJ  ; 
 ANI <=  RJI & TLN  |  RHI & TLN  |  ANI & tln  ; 
 ANJ <=  RJJ & TLN  |  RHJ & TLN  |  ANJ & tln  ; 
 RDI <=  IBI & TCC  |  IDI & TDC  |  IFI & TEC  |  IHI & TFC  ; 
 RHI <=  IBI & TCC  |  IDI & TDC  |  IFI & TEC  |  IHI & TFC  ; 
 qca <=  IJF  |  IJE  |  IJD  ; 
 qcb <=  IJF  |  IJE  |  ijd  ; 
 API <=  RJI & TLP  |  RHI & TLP  |  API & tlp  ; 
 APJ <=  RJJ & TLP  |  RHJ & TLP  |  APJ & tlp  ; 
 RDJ <=  IBJ & TCD  |  IDJ & TDD  |  IFJ & TED  |  IHJ & TFD  ; 
 RHJ <=  IBJ & TCD  |  IDJ & TDD  |  IFJ & TED  |  IHJ & TFD  ; 
 QDA <= IJA ; 
 QDB <= IJB ; 
 QDC <= IJC ; 
 CCC <=  BCC & JAK  |  BCC & JBK  ; 
 DCC <=  JAK & JAK  |  JBK & JBK  |  BCC  ; 
 CCD <=  BCD & JAL  |  BCD & JBL  ; 
 DCD <=  JAL & JAL  |  JBL & JBL  |  BCD  ; 
 kcc <=  gcc & hcc  |  GCC & HCC  |  tba  ; 
 kcg <=  gcg & hcc  |  GCG & HCC  |  tba  ; 
 kcd <=  gcd & hcd  |  GCD & HCD  |  tbb  ; 
 kch <=  gch & hcd  |  GCH & HCD  |  tbb  ; 
 kgd <=  ggd & hgd  |  GGD & HGD  |  tbd  ; 
 kgh <=  ggh & hgd  |  GGH & HGD  |  tbd  ; 
 kgc <=  ggc & hgc  |  GGC & HGC  |  tbc  ; 
 kgg <=  ggg & hgc  |  GGG & HGC  |  tbc  ; 
 CGC <=  BGC & JCK  |  BGC & JDK  ; 
 DGC <=  JCK & JCK  |  JDK & JDK  |  BGC  ; 
 CGD <=  BGD & JCL  |  BGD & JDL  ; 
 DGD <=  JCL & JCL  |  JDL & JDL  |  BGD  ; 
 BCC <=  jak & jbk & tia  |  JAK & TIA  |  JBK & TIC  ; 
 AAK <=  REK & TMA  |  RCK & TMA  |  AAK & tma  ; 
 AAL <=  REL & TMA  |  RCL & TMA  |  AAL & tma  ; 
 BCD <=  jal & jbl & tib  |  JAL & TIB  |  JBL & TID  ; 
 ACK <=  REK & TMC  |  RCK & TMC  |  ACK & tmc  ; 
 ACL <=  REL & TMC  |  RCL & TMC  |  ACL & tmc  ; 
 EAF <= qjb & QIA ; 
 EBF <= qjb & QIB ; 
 ECF <= qjb & QIC ; 
 EDF <= qjb & QID ; 
 RAK <=  KCC & pac  |  KCG & PAC  ; 
 RAL <=  KCD & pac  |  KCH & PAC  ; 
 AEK <=  REK & TME  |  RCK & TME  |  AEK & tme  ; 
 AEL <=  REL & TME  |  RCL & TME  |  AEL & tme  ; 
 QBA <= IKB ; 
 QBB <= QBA ; 
 QBC <= QBB ; 
 TLB <= FBB ; 
 TLJ <= FBB ; 
 TMB <= FBB ; 
 TMJ <= FBB ; 
 AGK <=  REK & TMG  |  RCK & TMG  |  AGK & tmg  ; 
 AGL <=  REL & TMG  |  RCL & TMG  |  AGL & tmg  ; 
 EEF <= qjd & QIE ; 
 EFF <= qjd & QIF ; 
 EGF <= qjd & QIG ; 
 EHF <= qjd & QIH ; 
 TLF <= FBF ; 
 TLN <= FBF ; 
 TMF <= FBF ; 
 TMN <= FBF ; 
 AIK <=  RFK & TLI  |  RDK & TLI  |  AIK & tli  ; 
 AIL <=  RFL & TLI  |  RDL & TLI  |  AIL & tli  ; 
 eif <= ZZI & QJB |  qia & qjb ; 
 ejf <= ZZI & QJB |  qib & qjb ; 
 ekf <= ZZI & QJB |  qic & qjb ; 
 RBK <=  KGC & pag  |  KGG & PAG  ; 
 RBL <=  KGD & pag  |  KGH & PAG  ; 
 AKK <=  RFK & TLK  |  RDK & TLK  |  AKK & tlk  ; 
 AKL <=  RFL & TLK  |  RDL & TLK  |  AKL & tlk  ; 
 elf <= ZZI & QJJ |  qid & qjj ; 
 epf <= ZZI & QJJ |  qih & qjj ; 
 BGC <=  jck & jdk & tie  |  JCK & TIE  |  JDK & TIG  ; 
 AMK <=  RFK & TLM  |  RDK & TLM  |  AMK & tlm  ; 
 AML <=  RFL & TLM  |  RDL & TLM  |  AML & tlm  ; 
 emf <= ZZI & QJD |  qie & qjd ; 
 enf <= ZZI & QJD |  qif & qjd ; 
 eof <= ZZI & QJD |  qig & qjd ; 
 BGD <=  jcl & jdl & tif  |  JCL & TIF  |  JDL & TIH  ; 
 AOK <=  RFK & TLO  |  RDK & TLO  |  AOK & tlo  ; 
 AOL <=  RFL & TLO  |  RDL & TLO  |  AOL & tlo  ; 
 ABK <=  RIK & TMB  |  RGK & TMB  |  ABK & tmb  ; 
 ABL <=  RIL & TMB  |  RGL & TMB  |  ABL & tmb  ; 
 RCK <=  IAK & TCA  |  ICK & TDA  |  IEK & TEA  |  IGK & TFA  ; 
 RGK <=  IAK & TCA  |  ICK & TDA  |  IEK & TEA  |  IGK & TFA  ; 
 qec <=  IIC  |  iib  |  IIA  ; 
 qed <=  IIC  |  iib  |  iia  ; 
 ADK <=  RIK & TMD  |  RGK & TMD  |  ADK & tmd  ; 
 ADL <=  RIL & TMD  |  RGL & TMD  |  ADL & tmd  ; 
 RCL <=  IAL & TCB  |  ICL & TDB  |  IEL & TEB  |  IGL & TFB  ; 
 RGL <=  IAL & TCB  |  ICL & TDB  |  IEL & TEB  |  IGL & TFB  ; 
 AFK <=  RIK & TMF  |  RGK & TMF  |  AFK & tmf  ; 
 AFL <=  RIL & TMF  |  RGL & TMF  |  AFL & tmf  ; 
 OGK <=  JEK  |  JFK  ; 
 SAK <=  JEK  |  JFK  ; 
 OAK <=  JEK  |  JFK  ; 
 OCK <=  JEK  |  JFK  ; 
 OEK <=  JEK  |  JFK  ; 
 AHK <=  RIK & TMH  |  RGK & TMH  |  AHK & tmh  ; 
 AHL <=  RIL & TMH  |  RGL & TMH  |  AHL & tmh  ; 
 OGL <=  JEL  |  JFL  ; 
 SAL <=  JEL  |  JFL  ; 
 OAL <=  JEL  |  JFL  ; 
 OCL <=  JEL  |  JFL  ; 
 OEL <=  JEL  |  JFL  ; 
 AJK <=  RJK & TLJ  |  RHK & TLJ  |  AJK & tlj  ; 
 AJL <=  RJL & TLJ  |  RHL & TLJ  |  AJL & tlj  ; 
 OHK <=  JGK  |  JHK  ; 
 SBK <=  JGK  |  JHK  ; 
 OBK <=  JGK  |  JHK  ; 
 ODK <=  JGK  |  JHK  ; 
 OFK <=  JGK  |  JHK  ; 
 ALK <=  RJK & TLL  |  RHK & TLL  |  ALK & tll  ; 
 ALL <=  RJL & TLL  |  RHL & TLL  |  ALL & tll  ; 
 OHL <=  JGL  |  JHL  ; 
 SBL <=  JGL  |  JHL  ; 
 OBL <=  JGL  |  JHL  ; 
 ODL <=  JGL  |  JHL  ; 
 OFL <=  JGL  |  JHL  ; 
 ANK <=  RJK & TLN  |  RHK & TLN  |  ANK & tln  ; 
 ANL <=  RJL & TLN  |  RHL & TLN  |  ANL & tln  ; 
 RDK <=  IBK & TCC  |  IDK & TDC  |  IFK & TEC  |  IHK & TFC  ; 
 RHK <=  IBK & TCC  |  IDK & TDC  |  IFK & TEC  |  IHK & TFC  ; 
 qcc <=  IJF  |  ije  |  IJD  ; 
 qcd <=  IJF  |  ije  |  ijd  ; 
 APK <=  RJK & TLP  |  RHK & TLP  |  APK & tlp  ; 
 APL <=  RJL & TLP  |  RHL & TLP  |  APL & tlp  ; 
 RDL <=  IBL & TCD  |  IDL & TDD  |  IFL & TED  |  IHL & TFD  ; 
 RHL <=  IBL & TCD  |  IDL & TDD  |  IFL & TED  |  IHL & TFD  ; 
 CDA <=  BDA & JAM  |  BDA & JBM  ; 
 DDA <=  JAM & JAM  |  JBM & JBM  |  BDA  ; 
 CDB <=  BDB & JAN  |  BDB & JBN  ; 
 DDB <=  JAN & JAN  |  JBN & JBN  |  BDB  ; 
 kda <=  hda  |  tba  ; 
 kde <=  HDA  |  tba  ; 
 kdb <=  gdb & hdb  |  GDB & HDB  |  tbb  ; 
 kdf <=  gdf & hdb  |  GDF & HDB  |  tbb  ; 
 QAE <= QAD ; 
 khb <=  ghb & hhb  |  GHB & HHB  |  tbd  ; 
 khf <=  ghf & hhb  |  GHF & HHB  |  tbd  ; 
 QAF <=  QAD & HAE & HBE & HCE & HDE  |  GAE & HBE & HCE & HDE  |  GBE & HCE & HDE  |  GCE & HDE & HDE  |  GDE  ; 
 kha <=  hha  |  tbc  ; 
 khe <=  HHA  |  tbc  ; 
 CHA <=  BHA & JCM  |  BHA & JDM  ; 
 DHA <=  JCM & JCM  |  JDM & JDM  |  BHA  ; 
 CHB <=  BHB & JCN  |  BHB & JDN  ; 
 DHB <=  JCN & JCN  |  JDN & JDN  |  BHB  ; 
 BDA <=  jam & jbm & tia  |  JAM & TIA  |  JBM & TIC  ; 
 AAM <=  REM & TMI  |  RCM & TMI  |  AAM & tmi  ; 
 AAN <=  REN & TMI  |  RCN & TMI  |  AAN & tmi  ; 
 BDB <=  jan & jbn & tib  |  JAN & TIB  |  JBN & TID  ; 
 ACM <=  REM & TMK  |  RCM & TMK  |  ACM & tmk  ; 
 ACN <=  REN & TMK  |  RCN & TMK  |  ACN & tmk  ; 
 EAG <= qja & QIA ; 
 EBG <= qja & QIB ; 
 ECG <= qja & QIC ; 
 EDG <= qja & QID ; 
 RAM <=  KDA & pad  |  KDE & PAD  ; 
 RAN <=  KDB & pad  |  KDF & PAD  ; 
 AEM <=  REM & TMM  |  RCM & TMM  |  AEM & tmm  ; 
 AEN <=  REN & TMM  |  RCN & TMM  |  AEN & tmm  ; 
 TLC <= FBC ; 
 TLK <= FBC ; 
 TMC <= FBC ; 
 TMK <= FBC ; 
 AGM <=  REM & TMO  |  RCM & TMO  |  AGM & tmo  ; 
 AGN <=  REN & TMO  |  RCN & TMO  |  AGN & tmo  ; 
 EEG <= qjc & QIE ; 
 EFG <= qjc & QIF ; 
 EGG <= qjc & QIG ; 
 EHG <= qjc & QIH ; 
 TLG <= FBG ; 
 TLO <= FBG ; 
 TMG <= FBG ; 
 TMO <= FBG ; 
 AIM <=  RFM & TLA  |  RDM & TLA  |  AIM & tla  ; 
 AIN <=  RFN & TLA  |  RDN & TLA  |  AIN & tla  ; 
 eig <= ZZI & QJA |  qia & qja ; 
 ejg <= ZZI & QJA |  qib & qja ; 
 ekg <= ZZI & QJA |  qic & qja ; 
 RBM <=  KHA & pah  |  KHE & PAH  ; 
 RBN <=  KHB & pah  |  KHF & PAH  ; 
 AKM <=  RFM & TLC  |  RDM & TLC  |  AKM & tlc  ; 
 AKN <=  RFN & TLC  |  RDN & TLC  |  AKN & tlc  ; 
 elg <= ZZI & QJK |  qid & qjk ; 
 epg <= ZZI & QJK |  qih & qjk ; 
 BHA <=  jcm & jdm & tie  |  JCM & TIE  |  JDM & TIG  ; 
 AMM <=  RFM & TLE  |  RDM & TLE  |  AMM & tle  ; 
 AMN <=  RFN & TLE  |  RDN & TLE  |  AMN & tle  ; 
 emg <= ZZI & QJC |  qie & qjc ; 
 eng <= ZZI & QJC |  qif & qjc ; 
 eog <= ZZI & QJC |  qig & qjc ; 
 BHB <=  jcn & jdn & tif  |  JCN & TIF  |  JDN & TIH  ; 
 AOM <=  RFM & TLG  |  RDM & TLG  |  AOM & tlg  ; 
 AON <=  RFN & TLG  |  RDN & TLG  |  AON & tlg  ; 
 ABM <=  RIM & TMJ  |  RGM & TMJ  |  ABM & tmj  ; 
 ABN <=  RIN & TMJ  |  RGN & TMJ  |  ABN & tmj  ; 
 RCM <=  IAM & TCA  |  ICM & TDA  |  IEM & TEA  |  IGM & TFA  ; 
 RGM <=  IAM & TCA  |  ICM & TDA  |  IEM & TEA  |  IGM & TFA  ; 
 qee <=  iic  |  IIB  |  IIA  ; 
 qef <=  iic  |  IIB  |  iia  ; 
 ADM <=  RIM & TML  |  RGM & TML  |  ADM & tml  ; 
 ADN <=  RIN & TML  |  RGN & TML  |  ADN & tml  ; 
 RCN <=  IAN & TCB  |  ICN & TDB  |  IEN & TEB  |  IGN & TFB  ; 
 RGN <=  IAN & TCB  |  ICN & TDB  |  IEN & TEB  |  IGN & TFB  ; 
 AFM <=  RIM & TMN  |  RGM & TMN  |  AFM & tmn  ; 
 AFN <=  RIN & TMN  |  RGN & TMN  |  AFN & tmn  ; 
 OGM <=  JEM  |  JFM  ; 
 SAM <=  JEM  |  JFM  ; 
 OAM <=  JEM  |  JFM  ; 
 OCM <=  JEM  |  JFM  ; 
 OEM <=  JEM  |  JFM  ; 
 AHM <=  RIM & TMP  |  RGM & TMP  |  AHM & tmp  ; 
 AHN <=  RIN & TMP  |  RGN & TMP  |  AHN & tmp  ; 
 OGN <=  JEN  |  JFN  ; 
 SAN <=  JEN  |  JFN  ; 
 OAN <=  JEN  |  JFN  ; 
 OCN <=  JEN  |  JFN  ; 
 OEN <=  JEN  |  JFN  ; 
 AJM <=  RJM & TLB  |  RHM & TLB  |  AJM & tlb  ; 
 AJN <=  RJN & TLB  |  RHN & TLB  |  AJN & tlb  ; 
 OHM <=  JGM  |  JHM  ; 
 SBM <=  JGM  |  JHM  ; 
 SCM <=  JGM  |  JHM  ; 
 OBM <=  JGM  |  JHM  ; 
 ODM <=  JGM  |  JHM  ; 
 OFM <=  JGM  |  JHM  ; 
 ALM <=  RJM & TLD  |  RHM & TLD  |  ALM & tld  ; 
 ALN <=  RJN & TLD  |  RHN & TLD  |  ALN & tld  ; 
 OHN <=  JGN  |  JHN  ; 
 SBN <=  JGN  |  JHN  ; 
 SCN <=  JGN  |  JHN  ; 
 OBN <=  JGN  |  JHN  ; 
 ODN <=  JGN  |  JHN  ; 
 OFN <=  JGN  |  JHN  ; 
 ANM <=  RJM & TLF  |  RHM & TLF  |  ANM & tlf  ; 
 ANN <=  RJN & TLF  |  RHN & TLF  |  ANN & tlf  ; 
 RDM <=  IBM & TCC  |  IDM & TDC  |  IFM & TEC  |  IHM & TFC  ; 
 RHM <=  IBM & TCC  |  IDM & TDC  |  IFM & TEC  |  IHM & TFC  ; 
 qce <=  ijf  |  IJE  |  IJD  ; 
 qcf <=  ijf  |  IJE  |  ijd  ; 
 APM <=  RJM & TLH  |  RHM & TLH  |  APM & tlh  ; 
 APN <=  RJN & TLH  |  RHN & TLH  |  APN & tlh  ; 
 RDN <=  IBN & TCD  |  IDN & TDD  |  IFN & TED  |  IHN & TFD  ; 
 RHN <=  IBN & TCD  |  IDN & TDD  |  IFN & TED  |  IHN & TFD  ; 
 CDC <=  BDC & JAO  |  BDC & JBO  ; 
 DDC <=  JAO & JAO  |  JBO & JBO  |  BDC  ; 
 CDD <=  BDD & JAP  |  BDD & JBP  ; 
 DDD <=  JAP & JAP  |  JBP & JBP  |  BDD  ; 
 kdc <=  gdc & hdc  |  GDC & HDC  |  tba  ; 
 kdg <=  gdg & hdc  |  GDG & HDC  |  tba  ; 
 kdd <=  gdd & hdd  |  GDD & HDD  |  tbb  ; 
 kdh <=  gdh & hdd  |  GDH & HDD  |  tbb  ; 
 khd <=  ghd & hhd  |  GHD & HHD  |  tbd  ; 
 khh <=  ghh & hhd  |  GHH & HHD  |  tbd  ; 
 khc <=  ghc & hhc  |  GHC & HHC  |  tbc  ; 
 khg <=  ghg & hhc  |  GHG & HHC  |  tbc  ; 
 CHC <=  BHC & JCO  |  BHC & JDO  ; 
 DHC <=  JCO & JCO  |  JDO & JDO  |  BHC  ; 
 CHD <=  BHD & JCP  |  BHD & JDP  ; 
 DHD <=  JCP & JCP  |  JDP & JDP  |  BHD  ; 
 BDC <=  jao & jbo & tia  |  JAO & TIA  |  JBO & TIC  ; 
 OMC <=  RIP & TMN  |  RGP & TMN  |  AFP & tmn  ; 
 AAO <=  REO & TMI  |  RCO & TMI  |  AAO & tmi  ; 
 AAP <=  REP & TMI  |  RCP & TMI  |  AAP & tmi  ; 
 BDD <=  jap & jbp & tib  |  JAP & TIB  |  JBP & TID  ; 
 OMD <=  RIP & TMP  |  RGP & TMP  |  AHP & tmp  ; 
 ACO <=  REO & TMK  |  RCO & TMK  |  ACO & tmk  ; 
 ACP <=  REP & TMK  |  RCP & TMK  |  ACP & tmk  ; 
 EAH <= qjb & QIA ; 
 EBH <= qjb & QIB ; 
 ECH <= qjb & QIC ; 
 EDH <= qjb & QID ; 
 RAO <=  KDC & pad  |  KDG & PAD  ; 
 RAP <=  KDD & pad  |  KDH & PAD  ; 
 AEO <=  REO & TMM  |  RCO & TMM  |  AEO & tmm  ; 
 AEP <=  REP & TMM  |  RCP & TMM  |  AEP & tmm  ; 
 TLD <= FBD ; 
 TLL <= FBD ; 
 TMD <= FBD ; 
 TML <= FBD ; 
 AGO <=  REO & TMO  |  RCO & TMO  |  AGO & tmo  ; 
 AGP <=  REP & TMO  |  RCP & TMO  |  AGP & tmo  ; 
 EEH <= qjd & QIE ; 
 EFH <= qjd & QIF ; 
 EGH <= qjd & QIG ; 
 EHH <= qjd & QIH ; 
 TLH <= FBH ; 
 TLP <= FBH ; 
 TMH <= FBH ; 
 TMP <= FBH ; 
 AIO <=  RFO & TLA  |  RDO & TLA  |  AIO & tla  ; 
 AIP <=  RFP & TLA  |  RDP & TLA  |  AIP & tla  ; 
 eih <= ZZI & QJB |  qia & qjb ; 
 ejh <= ZZI & QJB |  qib & qjb ; 
 ekh <= ZZI & QJB |  qic & qjb ; 
 RBO <=  KHC & pah  |  KHG & PAH  ; 
 RBP <=  KHD & pah  |  KHH & PAH  ; 
 AKO <=  RFO & TLC  |  RDO & TLC  |  AKO & tlc  ; 
 AKP <=  RFP & TLC  |  RDP & TLC  |  AKP & tlc  ; 
 elh <= ZZI & QJL |  qid & qjl ; 
 eph <= ZZI & QJL |  qih & qjl ; 
 BHC <=  jco & jdo & tie  |  JCO & TIE  |  JDO & TIG  ; 
 OMA <=  RIP & TMJ  |  RGP & TMJ  |  ABP & tmj  ; 
 AMO <=  RFO & TLE  |  RDO & TLE  |  AMO & tle  ; 
 AMP <=  RFP & TLE  |  RDP & TLE  |  AMP & tle  ; 
 emh <= ZZI & QJD |  qie & qjd ; 
 enh <= ZZI & QJD |  qif & qjd ; 
 eoh <= ZZI & QJD |  qig & qjd ; 
 BHD <=  jcp & jdp & tif  |  JCP & TIF  |  JDP & TIH  ; 
 OMB <=  RIP & TML  |  RGP & TML  |  ADP & tml  ; 
 AOO <=  RFO & TLG  |  RDO & TLG  |  AOO & tlg  ; 
 AOP <=  RFP & TLG  |  RDP & TLG  |  AOP & tlg  ; 
 ABO <=  RIO & TMJ  |  RGO & TMJ  |  ABO & tmj  ; 
 ABP <=  RIP & TMJ  |  RGP & TMJ  |  ABP & tmj  ; 
 RCO <=  IAO & TCA  |  ICO & TDA  |  IEO & TEA  |  IGO & TFA  ; 
 RGO <=  IAO & TCA  |  ICO & TDA  |  IEO & TEA  |  IGO & TFA  ; 
 qeg <=  iic  |  iib  |  IIA  ; 
 qeh <=  iic  |  iib  |  iia  ; 
 ADO <=  RIO & TML  |  RGO & TML  |  ADO & tml  ; 
 ADP <=  RIP & TML  |  RGP & TML  |  ADP & tml  ; 
 RCP <=  IAP & TCB  |  ICP & TDB  |  IEP & TEB  |  IGP & TFB  ; 
 RGP <=  IAP & TCB  |  ICP & TDB  |  IEP & TEB  |  IGP & TFB  ; 
 OKA <=  JIA  |  JIB  |  JIC  |  JID  ; 
 AFO <=  RIO & TMN  |  RGO & TMN  |  AFO & tmn  ; 
 AFP <=  RIP & TMN  |  RGP & TMN  |  AFP & tmn  ; 
 OGO <=  JEO  |  JFO  ; 
 SAO <=  JEO  |  JFO  ; 
 SCO <=  JEO  |  JFO  ; 
 OAO <=  JEO  |  JFO  ; 
 OCO <=  JEO  |  JFO  ; 
 OEO <=  JEO  |  JFO  ; 
 AHO <=  RIO & TMP  |  RGO & TMP  |  AHO & tmp  ; 
 AHP <=  RIP & TMP  |  RGP & TMP  |  AHP & tmp  ; 
 OGP <=  JEP  |  JFP  ; 
 SAP <=  JEP  |  JFP  ; 
 SCP <=  JEP  |  JFP  ; 
 OAP <=  JEP  |  JFP  ; 
 OCP <=  JEP  |  JFP  ; 
 OEP <=  JEP  |  JFP  ; 
 AJO <=  RJO & TLB  |  RHO & TLB  |  AJO & tlb  ; 
 AJP <=  RJP & TLB  |  RHP & TLB  |  AJP & tlb  ; 
 OHO <=  JGO  |  JHO  ; 
 SBO <=  JGO  |  JHO  ; 
 OBO <=  JGO  |  JHO  ; 
 ODO <=  JGO  |  JHO  ; 
 OFO <=  JGO  |  JHO  ; 
 ALO <=  RJO & TLD  |  RHO & TLD  |  ALO & tld  ; 
 ALP <=  RJP & TLD  |  RHP & TLD  |  ALP & tld  ; 
 OHP <=  JGP  |  JHP  ; 
 SBP <=  JGP  |  JHP  ; 
 OBP <=  JGP  |  JHP  ; 
 ODP <=  JGP  |  JHP  ; 
 OFP <=  JGP  |  JHP  ; 
 ANO <=  RJO & TLF  |  RHO & TLF  |  ANO & tlf  ; 
 ANP <=  RJP & TLF  |  RHP & TLF  |  ANP & tlf  ; 
 RDO <=  IBO & TCC  |  IDO & TDC  |  IFO & TEC  |  IHO & TFC  ; 
 RHO <=  IBO & TCC  |  IDO & TDC  |  IFO & TEC  |  IHO & TFC  ; 
 QKA <= IMA ; 
 ola <= sbp ; 
 APO <=  RJO & TLH  |  RHO & TLH  |  APO & tlh  ; 
 APP <=  RJP & TLH  |  RHP & TLH  |  APP & tlh  ; 
 RDP <=  IBP & TCD  |  IDP & TDD  |  IFP & TED  |  IHP & TFD  ; 
 RHP <=  IBP & TCD  |  IDP & TDD  |  IFP & TED  |  IHP & TFD  ; 
 OIJ <=  JIE  |  JIF  |  JIG  |  JIH  |  JIC  ; 
 OKB <=  JIE  |  JIF  |  JIG  |  JIH  |  JIC  ; 
 end 
end module
