module am( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFF, 
 IFG, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IHA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OIJ, 
 OIK, 
 OIL, 
 OIM, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OJM, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OLI, 
 OLJ, 
 OLK, 
 OLL, 
 OLM, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 OMG, 
 OMH, 
 OMI, 
 OMJ, 
 OMK, 
 OML, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ONG, 
 ONH, 
 ONI, 
 ONJ, 
 ONK, 
 ONL, 
 ONM, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OOG, 
 OOH, 
 OOI, 
 OOJ, 
 OOK, 
 OOL, 
 OOM, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPH, 
 OPI, 
 OPJ, 
 OPK, 
 OPL, 
OPM ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFF; 
 input IFG; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IHA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OIJ; 
 output OIK; 
 output OIL; 
 output OIM; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OJM; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OLI; 
 output OLJ; 
 output OLK; 
 output OLL; 
 output OLM; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output OMG; 
 output OMH; 
 output OMI; 
 output OMJ; 
 output OMK; 
 output OML; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ONG; 
 output ONH; 
 output ONI; 
 output ONJ; 
 output ONK; 
 output ONL; 
 output ONM; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OOG; 
 output OOH; 
 output OOI; 
 output OOJ; 
 output OOK; 
 output OOL; 
 output OOM; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPH; 
 output OPI; 
 output OPJ; 
 output OPK; 
 output OPL; 
 output OPM; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  AAQ ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ACQ ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  DGA ;
reg  DGC ;
reg  DGD ;
reg  dge ;
reg  DGF ;
reg  DGG ;
reg  dgh ;
reg  DGJ ;
reg  dgk ;
reg  DHA ;
reg  dhb ;
reg  DHC ;
reg  dhd ;
reg  DHE ;
reg  DHF ;
reg  DIA ;
reg  dib ;
reg  DIC ;
reg  did ;
reg  DIE ;
reg  dif ;
reg  DIG ;
reg  DJA ;
reg  djb ;
reg  DJC ;
reg  djd ;
reg  DJE ;
reg  djf ;
reg  DJG ;
reg  djh ;
reg  DKA ;
reg  dkb ;
reg  DKC ;
reg  dkd ;
reg  DKE ;
reg  dkf ;
reg  DKG ;
reg  dkh ;
reg  DKI ;
reg  DKJ ;
reg  DLA ;
reg  dlb ;
reg  DLC ;
reg  dld ;
reg  DLE ;
reg  dlf ;
reg  DLG ;
reg  dlh ;
reg  DLI ;
reg  dlj ;
reg  DLK ;
reg  DMA ;
reg  dmb ;
reg  DMC ;
reg  dmd ;
reg  DME ;
reg  dmf ;
reg  DMG ;
reg  dmh ;
reg  DMI ;
reg  dmj ;
reg  DMK ;
reg  dml ;
reg  DNA ;
reg  dnb ;
reg  DNC ;
reg  dnd ;
reg  DNE ;
reg  dnf ;
reg  DNG ;
reg  dnh ;
reg  DNI ;
reg  dnj ;
reg  DNK ;
reg  dnl ;
reg  DNM ;
reg  DNO ;
reg  DOA ;
reg  dob ;
reg  DOC ;
reg  dod ;
reg  DOE ;
reg  dof ;
reg  DOG ;
reg  doh ;
reg  DOI ;
reg  doj ;
reg  DOK ;
reg  dol ;
reg  DOM ;
reg  don ;
reg  DOO ;
reg  DPA ;
reg  dpb ;
reg  DPC ;
reg  dpd ;
reg  DPE ;
reg  dpf ;
reg  DPG ;
reg  dph ;
reg  DPI ;
reg  dpj ;
reg  DPK ;
reg  dpl ;
reg  DPM ;
reg  dpn ;
reg  DPO ;
reg  dpp ;
reg  DQA ;
reg  dqb ;
reg  DQC ;
reg  dqd ;
reg  DQE ;
reg  dqf ;
reg  DQG ;
reg  dqh ;
reg  DQI ;
reg  dqj ;
reg  DQK ;
reg  dql ;
reg  DQM ;
reg  dqn ;
reg  DQO ;
reg  dqp ;
reg  DQQ ;
reg  DQR ;
reg  DRA ;
reg  drb ;
reg  DRC ;
reg  drd ;
reg  DRE ;
reg  drf ;
reg  DRG ;
reg  drh ;
reg  DRI ;
reg  drj ;
reg  DRK ;
reg  drl ;
reg  DRM ;
reg  drn ;
reg  DRO ;
reg  drp ;
reg  DRQ ;
reg  drr ;
reg  DRS ;
reg  DSA ;
reg  dsb ;
reg  DSC ;
reg  dsd ;
reg  DSE ;
reg  dsf ;
reg  DSG ;
reg  dsh ;
reg  DSI ;
reg  dsj ;
reg  DSK ;
reg  dsl ;
reg  DSM ;
reg  dsn ;
reg  DSO ;
reg  dsp ;
reg  DSQ ;
reg  dsr ;
reg  DSS ;
reg  dst ;
reg  DTA ;
reg  dtb ;
reg  DTC ;
reg  dtd ;
reg  DTE ;
reg  dtf ;
reg  DTG ;
reg  dth ;
reg  DTI ;
reg  dtj ;
reg  DTK ;
reg  dtl ;
reg  DTM ;
reg  dtn ;
reg  DTO ;
reg  dtp ;
reg  DTQ ;
reg  dtr ;
reg  DTS ;
reg  dtt ;
reg  DTU ;
reg  DTV ;
reg  GAA ;
reg  gab ;
reg  GAC ;
reg  gad ;
reg  GAE ;
reg  GAF ;
reg  GBA ;
reg  gbb ;
reg  GBC ;
reg  gbd ;
reg  GBE ;
reg  GCA ;
reg  gcb ;
reg  GCC ;
reg  gcd ;
reg  GCE ;
reg  GDA ;
reg  gdb ;
reg  GDC ;
reg  gdd ;
reg  GDE ;
reg  GEA ;
reg  geb ;
reg  GEC ;
reg  ged ;
reg  GFA ;
reg  gfb ;
reg  GFC ;
reg  gfd ;
reg  GFE ;
reg  GGA ;
reg  ggb ;
reg  GGC ;
reg  ggd ;
reg  GHA ;
reg  ghb ;
reg  GHC ;
reg  ghd ;
reg  GHE ;
reg  GIA ;
reg  gib ;
reg  GIC ;
reg  gid ;
reg  GJA ;
reg  gjb ;
reg  GJC ;
reg  GJD ;
reg  GKA ;
reg  gkb ;
reg  GKC ;
reg  gkd ;
reg  GLA ;
reg  glb ;
reg  GLC ;
reg  GLD ;
reg  GMA ;
reg  gmb ;
reg  GMC ;
reg  GMD ;
reg  GNA ;
reg  gnb ;
reg  GNC ;
reg  GND ;
reg  GOA ;
reg  gob ;
reg  GOC ;
reg  GPA ;
reg  gpb ;
reg  GPC ;
reg  GQA ;
reg  gqb ;
reg  GQC ;
reg  GRA ;
reg  grb ;
reg  GRC ;
reg  GSA ;
reg  gsb ;
reg  GSC ;
reg  GTA ;
reg  gtb ;
reg  GUA ;
reg  gub ;
reg  GVA ;
reg  gvb ;
reg  GWA ;
reg  GWB ;
reg  GXA ;
reg  gxb ;
reg  GYA ;
reg  GYB ;
reg  GZA ;
reg  GZB ;
reg  GZD ;
reg  GZE ;
reg  GZF ;
reg  GZH ;
reg  GZK ;
reg  GZL ;
reg  GZM ;
reg  GZN ;
reg  JAA ;
reg  jab ;
reg  JAC ;
reg  JBA ;
reg  jbb ;
reg  JBC ;
reg  JCA ;
reg  jcb ;
reg  JCC ;
reg  JDA ;
reg  jdb ;
reg  JEA ;
reg  jeb ;
reg  JEC ;
reg  JFA ;
reg  jfb ;
reg  JGA ;
reg  jgb ;
reg  JGC ;
reg  JHA ;
reg  jhb ;
reg  JIA ;
reg  jib ;
reg  JJA ;
reg  jjb ;
reg  JKA ;
reg  jkb ;
reg  JLA ;
reg  jlb ;
reg  JMA ;
reg  jmb ;
reg  JNA ;
reg  JNB ;
reg  JOA ;
reg  JOB ;
reg  JPA ;
reg  JPB ;
reg  JQA ;
reg  JQB ;
reg  JRA ;
reg  JRB ;
reg  JSA ;
reg  JSB ;
reg  JTA ;
reg  JTB ;
reg  JUA ;
reg  JUB ;
reg  JVA ;
reg  JVB ;
reg  JWA ;
reg  JWB ;
reg  JXA ;
reg  JXB ;
reg  JYA ;
reg  JYB ;
reg  JZA ;
reg  JZC ;
reg  JZD ;
reg  JZE ;
reg  JZG ;
reg  JZI ;
reg  JZK ;
reg  JZL ;
reg  KBA ;
reg  kbb ;
reg  KBC ;
reg  KCA ;
reg  kcb ;
reg  KCC ;
reg  KDA ;
reg  kdb ;
reg  KDC ;
reg  KEA ;
reg  keb ;
reg  KFA ;
reg  kfb ;
reg  KFC ;
reg  KGA ;
reg  kgb ;
reg  KHA ;
reg  khb ;
reg  KHC ;
reg  KIA ;
reg  kib ;
reg  KJA ;
reg  kjb ;
reg  KKA ;
reg  kkb ;
reg  KLA ;
reg  klb ;
reg  KMA ;
reg  kmb ;
reg  KNA ;
reg  knb ;
reg  KOA ;
reg  KOB ;
reg  KPA ;
reg  KPB ;
reg  KQA ;
reg  KQB ;
reg  KRA ;
reg  KRB ;
reg  KSA ;
reg  KSB ;
reg  KTA ;
reg  KTB ;
reg  KUA ;
reg  KUB ;
reg  KVA ;
reg  KVB ;
reg  KWA ;
reg  KWB ;
reg  KXA ;
reg  KXB ;
reg  KYA ;
reg  KYB ;
reg  KZA ;
reg  KZB ;
reg  KZC ;
reg  KZE ;
reg  KZF ;
reg  KZG ;
reg  KZI ;
reg  KZJ ;
reg  KZL ;
reg  KZM ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  MAE ;
reg  MAF ;
reg  MAG ;
reg  MAH ;
reg  MAI ;
reg  MAJ ;
reg  MAK ;
reg  MAL ;
reg  MAM ;
reg  MAN ;
reg  MAO ;
reg  MAP ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  MBD ;
reg  MBE ;
reg  MBF ;
reg  MBG ;
reg  MBH ;
reg  MBI ;
reg  MBJ ;
reg  MBK ;
reg  MBL ;
reg  MBM ;
reg  MBN ;
reg  MBO ;
reg  MBP ;
reg  mca ;
reg  mcb ;
reg  mcc ;
reg  mcd ;
reg  mce ;
reg  mcf ;
reg  mcg ;
reg  mch ;
reg  mci ;
reg  mcj ;
reg  mck ;
reg  mcl ;
reg  mcm ;
reg  mcn ;
reg  mco ;
reg  mcp ;
reg  mda ;
reg  mdb ;
reg  mdc ;
reg  mdd ;
reg  mde ;
reg  mdf ;
reg  mdg ;
reg  mdh ;
reg  mdi ;
reg  MDJ ;
reg  MDK ;
reg  MDL ;
reg  MDM ;
reg  MDN ;
reg  MDQ ;
reg  MEA ;
reg  MEB ;
reg  MEC ;
reg  MED ;
reg  MEE ;
reg  MEF ;
reg  MEH ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  NBQ ;
reg  NEA ;
reg  NEB ;
reg  NEC ;
reg  NED ;
reg  nee ;
reg  nef ;
reg  neg ;
reg  NEH ;
reg  nei ;
reg  nej ;
reg  nek ;
reg  nel ;
reg  nem ;
reg  nen ;
reg  neo ;
reg  nep ;
reg  nfa ;
reg  nfb ;
reg  nfc ;
reg  nfd ;
reg  nfe ;
reg  nff ;
reg  nfg ;
reg  nfh ;
reg  nfi ;
reg  nfj ;
reg  nfk ;
reg  nfl ;
reg  nfm ;
reg  nfn ;
reg  nfo ;
reg  nfp ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  oia ;
reg  oib ;
reg  oic ;
reg  oid ;
reg  oie ;
reg  oif ;
reg  oig ;
reg  oih ;
reg  oii ;
reg  oij ;
reg  oik ;
reg  oil ;
reg  oim ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  OJK ;
reg  OJL ;
reg  OJM ;
reg  oka ;
reg  okb ;
reg  okc ;
reg  okd ;
reg  oke ;
reg  okf ;
reg  okg ;
reg  okh ;
reg  oki ;
reg  okj ;
reg  okk ;
reg  okl ;
reg  okm ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OLF ;
reg  OLG ;
reg  OLH ;
reg  OLI ;
reg  OLJ ;
reg  OLK ;
reg  OLL ;
reg  OLM ;
reg  oma ;
reg  omb ;
reg  omc ;
reg  omd ;
reg  ome ;
reg  omf ;
reg  omg ;
reg  omh ;
reg  omi ;
reg  omj ;
reg  omk ;
reg  oml ;
reg  omm ;
reg  ONA ;
reg  ONB ;
reg  ONC ;
reg  OND ;
reg  ONE ;
reg  ONF ;
reg  ONG ;
reg  ONH ;
reg  ONI ;
reg  ONJ ;
reg  ONK ;
reg  ONL ;
reg  ONM ;
reg  ooa ;
reg  oob ;
reg  ooc ;
reg  ood ;
reg  ooe ;
reg  oof ;
reg  oog ;
reg  ooh ;
reg  ooi ;
reg  ooj ;
reg  ook ;
reg  ool ;
reg  oom ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPH ;
reg  OPI ;
reg  OPJ ;
reg  OPK ;
reg  OPL ;
reg  OPM ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  pai ;
reg  pak ;
reg  PAL ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PCO ;
reg  PCP ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PDJ ;
reg  PDK ;
reg  PDL ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  PDP ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PEE ;
reg  PEF ;
reg  PEG ;
reg  PEH ;
reg  PEI ;
reg  PEJ ;
reg  PEK ;
reg  PEL ;
reg  PEM ;
reg  PEN ;
reg  PEO ;
reg  PEP ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PFE ;
reg  PFF ;
reg  PFG ;
reg  PFH ;
reg  PFI ;
reg  PFJ ;
reg  PFK ;
reg  PFL ;
reg  PFM ;
reg  PFN ;
reg  PFO ;
reg  PFP ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  PGD ;
reg  PGE ;
reg  PGF ;
reg  PGG ;
reg  PGH ;
reg  PGI ;
reg  PGJ ;
reg  PGK ;
reg  PGL ;
reg  PGM ;
reg  PGN ;
reg  PGO ;
reg  PGP ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aaq ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  acq ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  caa ;
wire  CAA ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  caf ;
wire  CAF ;
wire  cag ;
wire  CAG ;
wire  cah ;
wire  CAH ;
wire  cai ;
wire  CAI ;
wire  caj ;
wire  CAJ ;
wire  cak ;
wire  CAK ;
wire  cal ;
wire  CAL ;
wire  cam ;
wire  CAM ;
wire  can ;
wire  CAN ;
wire  cao ;
wire  CAO ;
wire  cap ;
wire  CAP ;
wire  cba ;
wire  CBA ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cbe ;
wire  CBE ;
wire  cbf ;
wire  CBF ;
wire  cbg ;
wire  CBG ;
wire  cbh ;
wire  CBH ;
wire  cbi ;
wire  CBI ;
wire  cbj ;
wire  CBJ ;
wire  cbk ;
wire  CBK ;
wire  cbl ;
wire  CBL ;
wire  cbm ;
wire  CBM ;
wire  cbn ;
wire  CBN ;
wire  cbo ;
wire  CBO ;
wire  cbp ;
wire  CBP ;
wire  cca ;
wire  CCA ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cce ;
wire  CCE ;
wire  ccf ;
wire  CCF ;
wire  ccg ;
wire  CCG ;
wire  cch ;
wire  CCH ;
wire  cci ;
wire  CCI ;
wire  ccj ;
wire  CCJ ;
wire  cck ;
wire  CCK ;
wire  ccl ;
wire  CCL ;
wire  ccm ;
wire  CCM ;
wire  ccn ;
wire  CCN ;
wire  cco ;
wire  CCO ;
wire  cda ;
wire  CDA ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cde ;
wire  CDE ;
wire  cdf ;
wire  CDF ;
wire  cdg ;
wire  CDG ;
wire  cdh ;
wire  CDH ;
wire  cdi ;
wire  CDI ;
wire  cdj ;
wire  CDJ ;
wire  cdk ;
wire  CDK ;
wire  cdl ;
wire  CDL ;
wire  cdm ;
wire  CDM ;
wire  cdn ;
wire  CDN ;
wire  cdo ;
wire  CDO ;
wire  cea ;
wire  CEA ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cee ;
wire  CEE ;
wire  cef ;
wire  CEF ;
wire  ceg ;
wire  CEG ;
wire  ceh ;
wire  CEH ;
wire  cei ;
wire  CEI ;
wire  cej ;
wire  CEJ ;
wire  cek ;
wire  CEK ;
wire  cel ;
wire  CEL ;
wire  cem ;
wire  CEM ;
wire  cen ;
wire  CEN ;
wire  cfa ;
wire  CFA ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cfe ;
wire  CFE ;
wire  cff ;
wire  CFF ;
wire  cfg ;
wire  CFG ;
wire  cfh ;
wire  CFH ;
wire  cfi ;
wire  CFI ;
wire  cfj ;
wire  CFJ ;
wire  cfk ;
wire  CFK ;
wire  cfl ;
wire  CFL ;
wire  cfm ;
wire  CFM ;
wire  cfn ;
wire  CFN ;
wire  cga ;
wire  CGA ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cge ;
wire  CGE ;
wire  cgf ;
wire  CGF ;
wire  cgg ;
wire  CGG ;
wire  cgh ;
wire  CGH ;
wire  cgi ;
wire  CGI ;
wire  cgj ;
wire  CGJ ;
wire  cgk ;
wire  CGK ;
wire  cgl ;
wire  CGL ;
wire  cgm ;
wire  CGM ;
wire  cha ;
wire  CHA ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  che ;
wire  CHE ;
wire  chf ;
wire  CHF ;
wire  chg ;
wire  CHG ;
wire  chh ;
wire  CHH ;
wire  chi ;
wire  CHI ;
wire  chj ;
wire  CHJ ;
wire  chk ;
wire  CHK ;
wire  chl ;
wire  CHL ;
wire  chm ;
wire  CHM ;
wire  cia ;
wire  CIA ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cie ;
wire  CIE ;
wire  cif ;
wire  CIF ;
wire  cig ;
wire  CIG ;
wire  cih ;
wire  CIH ;
wire  cii ;
wire  CII ;
wire  cij ;
wire  CIJ ;
wire  cik ;
wire  CIK ;
wire  cil ;
wire  CIL ;
wire  cja ;
wire  CJA ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cje ;
wire  CJE ;
wire  cjf ;
wire  CJF ;
wire  cjg ;
wire  CJG ;
wire  cjh ;
wire  CJH ;
wire  cji ;
wire  CJI ;
wire  cjj ;
wire  CJJ ;
wire  cjk ;
wire  CJK ;
wire  cjl ;
wire  CJL ;
wire  cka ;
wire  CKA ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cke ;
wire  CKE ;
wire  ckf ;
wire  CKF ;
wire  ckg ;
wire  CKG ;
wire  ckh ;
wire  CKH ;
wire  cki ;
wire  CKI ;
wire  ckj ;
wire  CKJ ;
wire  ckk ;
wire  CKK ;
wire  cla ;
wire  CLA ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cle ;
wire  CLE ;
wire  clf ;
wire  CLF ;
wire  clg ;
wire  CLG ;
wire  clh ;
wire  CLH ;
wire  cli ;
wire  CLI ;
wire  clj ;
wire  CLJ ;
wire  clk ;
wire  CLK ;
wire  cma ;
wire  CMA ;
wire  cmb ;
wire  CMB ;
wire  cmc ;
wire  CMC ;
wire  cmd ;
wire  CMD ;
wire  cme ;
wire  CME ;
wire  cmf ;
wire  CMF ;
wire  cmg ;
wire  CMG ;
wire  cmh ;
wire  CMH ;
wire  cmi ;
wire  CMI ;
wire  cmj ;
wire  CMJ ;
wire  cna ;
wire  CNA ;
wire  cnb ;
wire  CNB ;
wire  cnc ;
wire  CNC ;
wire  cnd ;
wire  CND ;
wire  cne ;
wire  CNE ;
wire  cnf ;
wire  CNF ;
wire  cng ;
wire  CNG ;
wire  cnh ;
wire  CNH ;
wire  cni ;
wire  CNI ;
wire  cnj ;
wire  CNJ ;
wire  coa ;
wire  COA ;
wire  cob ;
wire  COB ;
wire  coc ;
wire  COC ;
wire  cod ;
wire  COD ;
wire  coe ;
wire  COE ;
wire  cof ;
wire  COF ;
wire  cog ;
wire  COG ;
wire  coh ;
wire  COH ;
wire  coi ;
wire  COI ;
wire  cpa ;
wire  CPA ;
wire  cpb ;
wire  CPB ;
wire  cpc ;
wire  CPC ;
wire  cpd ;
wire  CPD ;
wire  cpe ;
wire  CPE ;
wire  cpf ;
wire  CPF ;
wire  cpg ;
wire  CPG ;
wire  cph ;
wire  CPH ;
wire  cpi ;
wire  CPI ;
wire  cqa ;
wire  CQA ;
wire  cqb ;
wire  CQB ;
wire  cqc ;
wire  CQC ;
wire  cqd ;
wire  CQD ;
wire  cqe ;
wire  CQE ;
wire  cqf ;
wire  CQF ;
wire  cqg ;
wire  CQG ;
wire  cqh ;
wire  CQH ;
wire  cra ;
wire  CRA ;
wire  crb ;
wire  CRB ;
wire  crc ;
wire  CRC ;
wire  crd ;
wire  CRD ;
wire  cre ;
wire  CRE ;
wire  crf ;
wire  CRF ;
wire  crg ;
wire  CRG ;
wire  crh ;
wire  CRH ;
wire  csa ;
wire  CSA ;
wire  csb ;
wire  CSB ;
wire  csc ;
wire  CSC ;
wire  csd ;
wire  CSD ;
wire  cse ;
wire  CSE ;
wire  csf ;
wire  CSF ;
wire  csg ;
wire  CSG ;
wire  cta ;
wire  CTA ;
wire  ctb ;
wire  CTB ;
wire  ctc ;
wire  CTC ;
wire  ctd ;
wire  CTD ;
wire  cte ;
wire  CTE ;
wire  ctf ;
wire  CTF ;
wire  ctg ;
wire  CTG ;
wire  cua ;
wire  CUA ;
wire  cub ;
wire  CUB ;
wire  cuc ;
wire  CUC ;
wire  cud ;
wire  CUD ;
wire  cue ;
wire  CUE ;
wire  cuf ;
wire  CUF ;
wire  cva ;
wire  CVA ;
wire  cvb ;
wire  CVB ;
wire  cvc ;
wire  CVC ;
wire  cvd ;
wire  CVD ;
wire  cve ;
wire  CVE ;
wire  cvf ;
wire  CVF ;
wire  cwa ;
wire  CWA ;
wire  cwb ;
wire  CWB ;
wire  cwc ;
wire  CWC ;
wire  cwd ;
wire  CWD ;
wire  cwe ;
wire  CWE ;
wire  cxa ;
wire  CXA ;
wire  cxb ;
wire  CXB ;
wire  cxc ;
wire  CXC ;
wire  cxd ;
wire  CXD ;
wire  cxe ;
wire  CXE ;
wire  cya ;
wire  CYA ;
wire  cyb ;
wire  CYB ;
wire  cyc ;
wire  CYC ;
wire  cyd ;
wire  CYD ;
wire  cza ;
wire  CZA ;
wire  czb ;
wire  CZB ;
wire  czc ;
wire  CZC ;
wire  czd ;
wire  CZD ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dca ;
wire  DCA ;
wire  dcb ;
wire  DCB ;
wire  dda ;
wire  DDA ;
wire  ddb ;
wire  DDB ;
wire  dea ;
wire  DEA ;
wire  dfa ;
wire  DFA ;
wire  dga ;
wire  dgc ;
wire  dgd ;
wire  DGE ;
wire  dgf ;
wire  dgg ;
wire  DGH ;
wire  dgj ;
wire  DGK ;
wire  dha ;
wire  DHB ;
wire  dhc ;
wire  DHD ;
wire  dhe ;
wire  dhf ;
wire  dia ;
wire  DIB ;
wire  dic ;
wire  DID ;
wire  die ;
wire  DIF ;
wire  dig ;
wire  dja ;
wire  DJB ;
wire  djc ;
wire  DJD ;
wire  dje ;
wire  DJF ;
wire  djg ;
wire  DJH ;
wire  dka ;
wire  DKB ;
wire  dkc ;
wire  DKD ;
wire  dke ;
wire  DKF ;
wire  dkg ;
wire  DKH ;
wire  dki ;
wire  dkj ;
wire  dla ;
wire  DLB ;
wire  dlc ;
wire  DLD ;
wire  dle ;
wire  DLF ;
wire  dlg ;
wire  DLH ;
wire  dli ;
wire  DLJ ;
wire  dlk ;
wire  dma ;
wire  DMB ;
wire  dmc ;
wire  DMD ;
wire  dme ;
wire  DMF ;
wire  dmg ;
wire  DMH ;
wire  dmi ;
wire  DMJ ;
wire  dmk ;
wire  DML ;
wire  dna ;
wire  DNB ;
wire  dnc ;
wire  DND ;
wire  dne ;
wire  DNF ;
wire  dng ;
wire  DNH ;
wire  dni ;
wire  DNJ ;
wire  dnk ;
wire  DNL ;
wire  dnm ;
wire  dno ;
wire  doa ;
wire  DOB ;
wire  doc ;
wire  DOD ;
wire  doe ;
wire  DOF ;
wire  dog ;
wire  DOH ;
wire  doi ;
wire  DOJ ;
wire  dok ;
wire  DOL ;
wire  dom ;
wire  DON ;
wire  doo ;
wire  dpa ;
wire  DPB ;
wire  dpc ;
wire  DPD ;
wire  dpe ;
wire  DPF ;
wire  dpg ;
wire  DPH ;
wire  dpi ;
wire  DPJ ;
wire  dpk ;
wire  DPL ;
wire  dpm ;
wire  DPN ;
wire  dpo ;
wire  DPP ;
wire  dqa ;
wire  DQB ;
wire  dqc ;
wire  DQD ;
wire  dqe ;
wire  DQF ;
wire  dqg ;
wire  DQH ;
wire  dqi ;
wire  DQJ ;
wire  dqk ;
wire  DQL ;
wire  dqm ;
wire  DQN ;
wire  dqo ;
wire  DQP ;
wire  dqq ;
wire  dqr ;
wire  dra ;
wire  DRB ;
wire  drc ;
wire  DRD ;
wire  dre ;
wire  DRF ;
wire  drg ;
wire  DRH ;
wire  dri ;
wire  DRJ ;
wire  drk ;
wire  DRL ;
wire  drm ;
wire  DRN ;
wire  dro ;
wire  DRP ;
wire  drq ;
wire  DRR ;
wire  drs ;
wire  dsa ;
wire  DSB ;
wire  dsc ;
wire  DSD ;
wire  dse ;
wire  DSF ;
wire  dsg ;
wire  DSH ;
wire  dsi ;
wire  DSJ ;
wire  dsk ;
wire  DSL ;
wire  dsm ;
wire  DSN ;
wire  dso ;
wire  DSP ;
wire  dsq ;
wire  DSR ;
wire  dss ;
wire  DST ;
wire  dta ;
wire  DTB ;
wire  dtc ;
wire  DTD ;
wire  dte ;
wire  DTF ;
wire  dtg ;
wire  DTH ;
wire  dti ;
wire  DTJ ;
wire  dtk ;
wire  DTL ;
wire  dtm ;
wire  DTN ;
wire  dto ;
wire  DTP ;
wire  dtq ;
wire  DTR ;
wire  dts ;
wire  DTT ;
wire  dtu ;
wire  dtv ;
wire  eaa ;
wire  EAA ;
wire  eba ;
wire  EBA ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  eda ;
wire  EDA ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eic ;
wire  EIC ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  ema ;
wire  EMA ;
wire  emb ;
wire  EMB ;
wire  emc ;
wire  EMC ;
wire  emd ;
wire  EMD ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  end ;
wire  END ;
wire  eoa ;
wire  EOA ;
wire  eob ;
wire  EOB ;
wire  eoc ;
wire  EOC ;
wire  eod ;
wire  EOD ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  eqa ;
wire  EQA ;
wire  eqb ;
wire  EQB ;
wire  eqc ;
wire  EQC ;
wire  eqd ;
wire  EQD ;
wire  era ;
wire  ERA ;
wire  erb ;
wire  ERB ;
wire  erc ;
wire  ERC ;
wire  erd ;
wire  ERD ;
wire  esa ;
wire  ESA ;
wire  esb ;
wire  ESB ;
wire  esc ;
wire  ESC ;
wire  esd ;
wire  ESD ;
wire  ese ;
wire  ESE ;
wire  eta ;
wire  ETA ;
wire  etb ;
wire  ETB ;
wire  etc ;
wire  ETC ;
wire  etd ;
wire  ETD ;
wire  ete ;
wire  ETE ;
wire  eua ;
wire  EUA ;
wire  eub ;
wire  EUB ;
wire  euc ;
wire  EUC ;
wire  eud ;
wire  EUD ;
wire  eue ;
wire  EUE ;
wire  euf ;
wire  EUF ;
wire  eva ;
wire  EVA ;
wire  evb ;
wire  EVB ;
wire  evc ;
wire  EVC ;
wire  evd ;
wire  EVD ;
wire  eve ;
wire  EVE ;
wire  ewa ;
wire  EWA ;
wire  ewb ;
wire  EWB ;
wire  ewc ;
wire  EWC ;
wire  ewd ;
wire  EWD ;
wire  ewe ;
wire  EWE ;
wire  ewf ;
wire  EWF ;
wire  exa ;
wire  EXA ;
wire  exb ;
wire  EXB ;
wire  exc ;
wire  EXC ;
wire  exd ;
wire  EXD ;
wire  exe ;
wire  EXE ;
wire  exf ;
wire  EXF ;
wire  eya ;
wire  EYA ;
wire  eyb ;
wire  EYB ;
wire  eyc ;
wire  EYC ;
wire  eyd ;
wire  EYD ;
wire  eye ;
wire  EYE ;
wire  eyf ;
wire  EYF ;
wire  eyg ;
wire  EYG ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fea ;
wire  FEA ;
wire  feb ;
wire  FEB ;
wire  fec ;
wire  FEC ;
wire  fed ;
wire  FED ;
wire  fee ;
wire  FEE ;
wire  fef ;
wire  FEF ;
wire  feg ;
wire  FEG ;
wire  ffa ;
wire  FFA ;
wire  ffb ;
wire  FFB ;
wire  ffc ;
wire  FFC ;
wire  ffd ;
wire  FFD ;
wire  ffe ;
wire  FFE ;
wire  fff ;
wire  FFF ;
wire  ffg ;
wire  FFG ;
wire  ffh ;
wire  FFH ;
wire  fga ;
wire  FGA ;
wire  fgb ;
wire  FGB ;
wire  fgc ;
wire  FGC ;
wire  fgd ;
wire  FGD ;
wire  fge ;
wire  FGE ;
wire  fgf ;
wire  FGF ;
wire  fgg ;
wire  FGG ;
wire  fgh ;
wire  FGH ;
wire  gaa ;
wire  GAB ;
wire  gac ;
wire  GAD ;
wire  gae ;
wire  gaf ;
wire  gba ;
wire  GBB ;
wire  gbc ;
wire  GBD ;
wire  gbe ;
wire  gca ;
wire  GCB ;
wire  gcc ;
wire  GCD ;
wire  gce ;
wire  gda ;
wire  GDB ;
wire  gdc ;
wire  GDD ;
wire  gde ;
wire  gea ;
wire  GEB ;
wire  gec ;
wire  GED ;
wire  gfa ;
wire  GFB ;
wire  gfc ;
wire  GFD ;
wire  gfe ;
wire  gga ;
wire  GGB ;
wire  ggc ;
wire  GGD ;
wire  gha ;
wire  GHB ;
wire  ghc ;
wire  GHD ;
wire  ghe ;
wire  gia ;
wire  GIB ;
wire  gic ;
wire  GID ;
wire  gja ;
wire  GJB ;
wire  gjc ;
wire  gjd ;
wire  gka ;
wire  GKB ;
wire  gkc ;
wire  GKD ;
wire  gla ;
wire  GLB ;
wire  glc ;
wire  gld ;
wire  gma ;
wire  GMB ;
wire  gmc ;
wire  gmd ;
wire  gna ;
wire  GNB ;
wire  gnc ;
wire  gnd ;
wire  goa ;
wire  GOB ;
wire  goc ;
wire  gpa ;
wire  GPB ;
wire  gpc ;
wire  gqa ;
wire  GQB ;
wire  gqc ;
wire  gra ;
wire  GRB ;
wire  grc ;
wire  gsa ;
wire  GSB ;
wire  gsc ;
wire  gta ;
wire  GTB ;
wire  gua ;
wire  GUB ;
wire  gva ;
wire  GVB ;
wire  gwa ;
wire  gwb ;
wire  gxa ;
wire  GXB ;
wire  gya ;
wire  gyb ;
wire  gza ;
wire  gzb ;
wire  gzd ;
wire  gze ;
wire  gzf ;
wire  gzh ;
wire  gzk ;
wire  gzl ;
wire  gzm ;
wire  gzn ;
wire  haa ;
wire  HAA ;
wire  hab ;
wire  HAB ;
wire  hac ;
wire  HAC ;
wire  had ;
wire  HAD ;
wire  hba ;
wire  HBA ;
wire  hbb ;
wire  HBB ;
wire  hbc ;
wire  HBC ;
wire  hbd ;
wire  HBD ;
wire  hca ;
wire  HCA ;
wire  hcb ;
wire  HCB ;
wire  hcd ;
wire  HCD ;
wire  hce ;
wire  HCE ;
wire  hda ;
wire  HDA ;
wire  hdb ;
wire  HDB ;
wire  hdc ;
wire  HDC ;
wire  hdd ;
wire  HDD ;
wire  hea ;
wire  HEA ;
wire  heb ;
wire  HEB ;
wire  hec ;
wire  HEC ;
wire  hfa ;
wire  HFA ;
wire  hfb ;
wire  HFB ;
wire  hfc ;
wire  HFC ;
wire  hfd ;
wire  HFD ;
wire  hga ;
wire  HGA ;
wire  hgb ;
wire  HGB ;
wire  hgc ;
wire  HGC ;
wire  hha ;
wire  HHA ;
wire  hhb ;
wire  HHB ;
wire  hhc ;
wire  HHC ;
wire  hhd ;
wire  HHD ;
wire  hia ;
wire  HIA ;
wire  hib ;
wire  HIB ;
wire  hic ;
wire  HIC ;
wire  hja ;
wire  HJA ;
wire  hjb ;
wire  HJB ;
wire  hjc ;
wire  HJC ;
wire  hka ;
wire  HKA ;
wire  hkb ;
wire  HKB ;
wire  hkc ;
wire  HKC ;
wire  hla ;
wire  HLA ;
wire  hlb ;
wire  HLB ;
wire  hlc ;
wire  HLC ;
wire  hma ;
wire  HMA ;
wire  hmb ;
wire  HMB ;
wire  hmc ;
wire  HMC ;
wire  hna ;
wire  HNA ;
wire  hnb ;
wire  HNB ;
wire  hoa ;
wire  HOA ;
wire  hob ;
wire  HOB ;
wire  hpa ;
wire  HPA ;
wire  hpb ;
wire  HPB ;
wire  hqa ;
wire  HQA ;
wire  hqb ;
wire  HQB ;
wire  hra ;
wire  HRA ;
wire  hrb ;
wire  HRB ;
wire  hsa ;
wire  HSA ;
wire  hsb ;
wire  HSB ;
wire  hta ;
wire  HTA ;
wire  htb ;
wire  HTB ;
wire  hua ;
wire  HUA ;
wire  hub ;
wire  HUB ;
wire  hva ;
wire  HVA ;
wire  hvb ;
wire  HVB ;
wire  hwa ;
wire  HWA ;
wire  hwb ;
wire  HWB ;
wire  hxa ;
wire  HXA ;
wire  hxb ;
wire  HXB ;
wire  hya ;
wire  HYA ;
wire  hyb ;
wire  HYB ;
wire  hza ;
wire  HZA ;
wire  hzb ;
wire  HZB ;
wire  hzc ;
wire  HZC ;
wire  hze ;
wire  HZE ;
wire  hzf ;
wire  HZF ;
wire  hzg ;
wire  HZG ;
wire  hzi ;
wire  HZI ;
wire  hzk ;
wire  HZK ;
wire  hzl ;
wire  HZL ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iff ;
wire  ifg ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  iha ;
wire  jaa ;
wire  JAB ;
wire  jac ;
wire  jba ;
wire  JBB ;
wire  jbc ;
wire  jca ;
wire  JCB ;
wire  jcc ;
wire  jda ;
wire  JDB ;
wire  jea ;
wire  JEB ;
wire  jec ;
wire  jfa ;
wire  JFB ;
wire  jga ;
wire  JGB ;
wire  jgc ;
wire  jha ;
wire  JHB ;
wire  jia ;
wire  JIB ;
wire  jja ;
wire  JJB ;
wire  jka ;
wire  JKB ;
wire  jla ;
wire  JLB ;
wire  jma ;
wire  JMB ;
wire  jna ;
wire  jnb ;
wire  joa ;
wire  job ;
wire  jpa ;
wire  jpb ;
wire  jqa ;
wire  jqb ;
wire  jra ;
wire  jrb ;
wire  jsa ;
wire  jsb ;
wire  jta ;
wire  jtb ;
wire  jua ;
wire  jub ;
wire  jva ;
wire  jvb ;
wire  jwa ;
wire  jwb ;
wire  jxa ;
wire  jxb ;
wire  jya ;
wire  jyb ;
wire  jza ;
wire  jzc ;
wire  jzd ;
wire  jze ;
wire  jzg ;
wire  jzi ;
wire  jzk ;
wire  jzl ;
wire  kba ;
wire  KBB ;
wire  kbc ;
wire  kca ;
wire  KCB ;
wire  kcc ;
wire  kda ;
wire  KDB ;
wire  kdc ;
wire  kea ;
wire  KEB ;
wire  kfa ;
wire  KFB ;
wire  kfc ;
wire  kga ;
wire  KGB ;
wire  kha ;
wire  KHB ;
wire  khc ;
wire  kia ;
wire  KIB ;
wire  kja ;
wire  KJB ;
wire  kka ;
wire  KKB ;
wire  kla ;
wire  KLB ;
wire  kma ;
wire  KMB ;
wire  kna ;
wire  KNB ;
wire  koa ;
wire  kob ;
wire  kpa ;
wire  kpb ;
wire  kqa ;
wire  kqb ;
wire  kra ;
wire  krb ;
wire  ksa ;
wire  ksb ;
wire  kta ;
wire  ktb ;
wire  kua ;
wire  kub ;
wire  kva ;
wire  kvb ;
wire  kwa ;
wire  kwb ;
wire  kxa ;
wire  kxb ;
wire  kya ;
wire  kyb ;
wire  kza ;
wire  kzb ;
wire  kzc ;
wire  kze ;
wire  kzf ;
wire  kzg ;
wire  kzi ;
wire  kzj ;
wire  kzl ;
wire  kzm ;
wire  lba ;
wire  LBA ;
wire  lbb ;
wire  LBB ;
wire  lbc ;
wire  LBC ;
wire  lbd ;
wire  LBD ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lcc ;
wire  LCC ;
wire  lcd ;
wire  LCD ;
wire  lce ;
wire  LCE ;
wire  lda ;
wire  LDA ;
wire  ldb ;
wire  LDB ;
wire  ldc ;
wire  LDC ;
wire  ldd ;
wire  LDD ;
wire  lea ;
wire  LEA ;
wire  leb ;
wire  LEB ;
wire  lec ;
wire  LEC ;
wire  led ;
wire  LED ;
wire  lfa ;
wire  LFA ;
wire  lfb ;
wire  LFB ;
wire  lfc ;
wire  LFC ;
wire  lfd ;
wire  LFD ;
wire  lga ;
wire  LGA ;
wire  lgb ;
wire  LGB ;
wire  lgc ;
wire  LGC ;
wire  lgd ;
wire  LGD ;
wire  lha ;
wire  LHA ;
wire  lhb ;
wire  LHB ;
wire  lhc ;
wire  LHC ;
wire  lhd ;
wire  LHD ;
wire  lia ;
wire  LIA ;
wire  lib ;
wire  LIB ;
wire  lic ;
wire  LIC ;
wire  lja ;
wire  LJA ;
wire  ljb ;
wire  LJB ;
wire  ljc ;
wire  LJC ;
wire  lka ;
wire  LKA ;
wire  lkb ;
wire  LKB ;
wire  lkc ;
wire  LKC ;
wire  lla ;
wire  LLA ;
wire  llb ;
wire  LLB ;
wire  llc ;
wire  LLC ;
wire  lma ;
wire  LMA ;
wire  lmb ;
wire  LMB ;
wire  lmc ;
wire  LMC ;
wire  lna ;
wire  LNA ;
wire  lnb ;
wire  LNB ;
wire  lnc ;
wire  LNC ;
wire  loa ;
wire  LOA ;
wire  lob ;
wire  LOB ;
wire  loc ;
wire  LOC ;
wire  lpa ;
wire  LPA ;
wire  lpb ;
wire  LPB ;
wire  lpc ;
wire  LPC ;
wire  lqa ;
wire  LQA ;
wire  lqb ;
wire  LQB ;
wire  lqc ;
wire  LQC ;
wire  lra ;
wire  LRA ;
wire  lrb ;
wire  LRB ;
wire  lrc ;
wire  LRC ;
wire  lsa ;
wire  LSA ;
wire  lsb ;
wire  LSB ;
wire  lsc ;
wire  LSC ;
wire  lta ;
wire  LTA ;
wire  ltb ;
wire  LTB ;
wire  ltc ;
wire  LTC ;
wire  lua ;
wire  LUA ;
wire  lub ;
wire  LUB ;
wire  luc ;
wire  LUC ;
wire  lva ;
wire  LVA ;
wire  lvb ;
wire  LVB ;
wire  lvc ;
wire  LVC ;
wire  lwa ;
wire  LWA ;
wire  lwb ;
wire  LWB ;
wire  lwc ;
wire  LWC ;
wire  lxa ;
wire  LXA ;
wire  lxb ;
wire  LXB ;
wire  lxc ;
wire  LXC ;
wire  lya ;
wire  LYA ;
wire  lyb ;
wire  LYB ;
wire  lyc ;
wire  LYC ;
wire  lza ;
wire  LZA ;
wire  lzb ;
wire  LZB ;
wire  lzc ;
wire  LZC ;
wire  lzd ;
wire  LZD ;
wire  lze ;
wire  LZE ;
wire  lzf ;
wire  LZF ;
wire  lzg ;
wire  LZG ;
wire  lzh ;
wire  LZH ;
wire  lzi ;
wire  LZI ;
wire  lzj ;
wire  LZJ ;
wire  lzk ;
wire  LZK ;
wire  lzl ;
wire  LZL ;
wire  lzm ;
wire  LZM ;
wire  lzn ;
wire  LZN ;
wire  lzo ;
wire  LZO ;
wire  lzp ;
wire  LZP ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  mae ;
wire  maf ;
wire  mag ;
wire  mah ;
wire  mai ;
wire  maj ;
wire  mak ;
wire  mal ;
wire  mam ;
wire  man ;
wire  mao ;
wire  map ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  mbd ;
wire  mbe ;
wire  mbf ;
wire  mbg ;
wire  mbh ;
wire  mbi ;
wire  mbj ;
wire  mbk ;
wire  mbl ;
wire  mbm ;
wire  mbn ;
wire  mbo ;
wire  mbp ;
wire  MCA ;
wire  MCB ;
wire  MCC ;
wire  MCD ;
wire  MCE ;
wire  MCF ;
wire  MCG ;
wire  MCH ;
wire  MCI ;
wire  MCJ ;
wire  MCK ;
wire  MCL ;
wire  MCM ;
wire  MCN ;
wire  MCO ;
wire  MCP ;
wire  MDA ;
wire  MDB ;
wire  MDC ;
wire  MDD ;
wire  MDE ;
wire  MDF ;
wire  MDG ;
wire  MDH ;
wire  MDI ;
wire  mdj ;
wire  mdk ;
wire  mdl ;
wire  mdm ;
wire  mdn ;
wire  mdq ;
wire  mea ;
wire  meb ;
wire  mec ;
wire  med ;
wire  mee ;
wire  mef ;
wire  meh ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  nbq ;
wire  nea ;
wire  neb ;
wire  nec ;
wire  ned ;
wire  NEE ;
wire  NEF ;
wire  NEG ;
wire  neh ;
wire  NEI ;
wire  NEJ ;
wire  NEK ;
wire  NEL ;
wire  NEM ;
wire  NEN ;
wire  NEO ;
wire  NEP ;
wire  NFA ;
wire  NFB ;
wire  NFC ;
wire  NFD ;
wire  NFE ;
wire  NFF ;
wire  NFG ;
wire  NFH ;
wire  NFI ;
wire  NFJ ;
wire  NFK ;
wire  NFL ;
wire  NFM ;
wire  NFN ;
wire  NFO ;
wire  NFP ;
wire  nhb ;
wire  NHB ;
wire  nhc ;
wire  NHC ;
wire  nhd ;
wire  NHD ;
wire  nhe ;
wire  NHE ;
wire  nib ;
wire  NIB ;
wire  nic ;
wire  NIC ;
wire  nid ;
wire  NID ;
wire  nie ;
wire  NIE ;
wire  njb ;
wire  NJB ;
wire  njc ;
wire  NJC ;
wire  njd ;
wire  NJD ;
wire  nje ;
wire  NJE ;
wire  nkb ;
wire  NKB ;
wire  nkc ;
wire  NKC ;
wire  nkd ;
wire  NKD ;
wire  nke ;
wire  NKE ;
wire  nlb ;
wire  NLB ;
wire  nlc ;
wire  NLC ;
wire  nld ;
wire  NLD ;
wire  nle ;
wire  NLE ;
wire  nmb ;
wire  NMB ;
wire  nmc ;
wire  NMC ;
wire  nmd ;
wire  NMD ;
wire  nme ;
wire  NME ;
wire  nnb ;
wire  NNB ;
wire  nnc ;
wire  NNC ;
wire  nnd ;
wire  NND ;
wire  nne ;
wire  NNE ;
wire  npb ;
wire  NPB ;
wire  npc ;
wire  NPC ;
wire  npd ;
wire  NPD ;
wire  nqb ;
wire  NQB ;
wire  nqc ;
wire  NQC ;
wire  nqd ;
wire  NQD ;
wire  nrb ;
wire  NRB ;
wire  nrc ;
wire  NRC ;
wire  nrd ;
wire  NRD ;
wire  nsb ;
wire  NSB ;
wire  nsc ;
wire  NSC ;
wire  nsd ;
wire  NSD ;
wire  ntb ;
wire  NTB ;
wire  ntc ;
wire  NTC ;
wire  ntd ;
wire  NTD ;
wire  nub ;
wire  NUB ;
wire  nuc ;
wire  NUC ;
wire  nud ;
wire  NUD ;
wire  nvb ;
wire  NVB ;
wire  nvc ;
wire  NVC ;
wire  nvd ;
wire  NVD ;
wire  nxb ;
wire  NXB ;
wire  nxc ;
wire  NXC ;
wire  nxd ;
wire  NXD ;
wire  nxe ;
wire  NXE ;
wire  nxf ;
wire  NXF ;
wire  nxg ;
wire  NXG ;
wire  nxi ;
wire  NXI ;
wire  nxj ;
wire  NXJ ;
wire  nxk ;
wire  NXK ;
wire  nxl ;
wire  NXL ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OIA ;
wire  OIB ;
wire  OIC ;
wire  OID ;
wire  OIE ;
wire  OIF ;
wire  OIG ;
wire  OIH ;
wire  OII ;
wire  OIJ ;
wire  OIK ;
wire  OIL ;
wire  OIM ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  ojk ;
wire  ojl ;
wire  ojm ;
wire  OKA ;
wire  OKB ;
wire  OKC ;
wire  OKD ;
wire  OKE ;
wire  OKF ;
wire  OKG ;
wire  OKH ;
wire  OKI ;
wire  OKJ ;
wire  OKK ;
wire  OKL ;
wire  OKM ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  olf ;
wire  olg ;
wire  olh ;
wire  oli ;
wire  olj ;
wire  olk ;
wire  oll ;
wire  olm ;
wire  OMA ;
wire  OMB ;
wire  OMC ;
wire  OMD ;
wire  OME ;
wire  OMF ;
wire  OMG ;
wire  OMH ;
wire  OMI ;
wire  OMJ ;
wire  OMK ;
wire  OML ;
wire  OMM ;
wire  ona ;
wire  onb ;
wire  onc ;
wire  ond ;
wire  one ;
wire  onf ;
wire  ong ;
wire  onh ;
wire  oni ;
wire  onj ;
wire  onk ;
wire  onl ;
wire  onm ;
wire  OOA ;
wire  OOB ;
wire  OOC ;
wire  OOD ;
wire  OOE ;
wire  OOF ;
wire  OOG ;
wire  OOH ;
wire  OOI ;
wire  OOJ ;
wire  OOK ;
wire  OOL ;
wire  OOM ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  oph ;
wire  opi ;
wire  opj ;
wire  opk ;
wire  opl ;
wire  opm ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  PAI ;
wire  PAK ;
wire  pal ;
wire  pam ;
wire  PAM ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pco ;
wire  pcp ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pdj ;
wire  pdk ;
wire  pdl ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  pdp ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pee ;
wire  pef ;
wire  peg ;
wire  peh ;
wire  pei ;
wire  pej ;
wire  pek ;
wire  pel ;
wire  pem ;
wire  pen ;
wire  peo ;
wire  pep ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pfe ;
wire  pff ;
wire  pfg ;
wire  pfh ;
wire  pfi ;
wire  pfj ;
wire  pfk ;
wire  pfl ;
wire  pfm ;
wire  pfn ;
wire  pfo ;
wire  pfp ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  pgd ;
wire  pge ;
wire  pgf ;
wire  pgg ;
wire  pgh ;
wire  pgi ;
wire  pgj ;
wire  pgk ;
wire  pgl ;
wire  pgm ;
wire  pgn ;
wire  pgo ;
wire  pgp ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  teg ;
wire  TEG ;
wire  teh ;
wire  TEH ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign aal = ~AAL;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign man = ~MAN;  //complement 
assign MCN = ~mcn;  //complement 
assign drq = ~DRQ;  //complement 
assign DRR = ~drr;  //complement 
assign nea = ~NEA;  //complement 
assign neb = ~NEB;  //complement 
assign nec = ~NEC;  //complement 
assign mdm = ~MDM;  //complement 
assign ojg = ~OJG;  //complement 
assign olg = ~OLG;  //complement 
assign ong = ~ONG;  //complement 
assign opg = ~OPG;  //complement 
assign mao = ~MAO;  //complement 
assign MCO = ~mco;  //complement 
assign dsa = ~DSA;  //complement 
assign DSB = ~dsb;  //complement 
assign dga = ~DGA;  //complement 
assign dgc = ~DGC;  //complement 
assign map = ~MAP;  //complement 
assign MCP = ~mcp;  //complement 
assign dsc = ~DSC;  //complement 
assign DSD = ~dsd;  //complement 
assign dnm = ~DNM;  //complement 
assign dno = ~DNO;  //complement 
assign mba = ~MBA;  //complement 
assign MDA = ~mda;  //complement 
assign dse = ~DSE;  //complement 
assign DSF = ~dsf;  //complement 
assign dqr = ~DQR;  //complement 
assign gzn = ~GZN;  //complement 
assign mbb = ~MBB;  //complement 
assign MDB = ~mdb;  //complement 
assign mdq = ~MDQ;  //complement 
assign dsg = ~DSG;  //complement 
assign DSH = ~dsh;  //complement 
assign gjd = ~GJD;  //complement 
assign ned = ~NED;  //complement 
assign mbc = ~MBC;  //complement 
assign MDC = ~mdc;  //complement 
assign dsi = ~DSI;  //complement 
assign DSJ = ~dsj;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign mbd = ~MBD;  //complement 
assign MDD = ~mdd;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign aak = ~AAK;  //complement 
assign mbe = ~MBE;  //complement 
assign MDE = ~mde;  //complement 
assign dsk = ~DSK;  //complement 
assign DSL = ~dsl;  //complement 
assign dsm = ~DSM;  //complement 
assign DSN = ~dsn;  //complement 
assign dgd = ~DGD;  //complement 
assign DGE = ~dge;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign FGA =  DTB & dtd & dtf  |  dtb & DTD & dtf  |  dtb & dtd & DTF  |  DTB & DTD & DTF  ; 
assign fga = ~FGA; //complement 
assign fgb =  DTB & dtd & dtf  |  dtb & DTD & dtf  |  dtb & dtd & DTF  |  dtb & dtd & dtf  ; 
assign FGB = ~fgb;  //complement 
assign FGC =  DTH & dtj & dtl  |  dth & DTJ & dtl  |  dth & dtj & DTL  |  DTH & DTJ & DTL  ; 
assign fgc = ~FGC; //complement 
assign fgd =  DTH & dtj & dtl  |  dth & DTJ & dtl  |  dth & dtj & DTL  |  dth & dtj & dtl  ; 
assign FGD = ~fgd;  //complement 
assign dgg = ~DGG;  //complement 
assign DGH = ~dgh;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign abk = ~ABK;  //complement 
assign FGE =  DTN & dtp & dtr  |  dtn & DTP & dtr  |  dtn & dtp & DTR  |  DTN & DTP & DTR  ; 
assign fge = ~FGE; //complement 
assign fgf =  DTN & dtp & dtr  |  dtn & DTP & dtr  |  dtn & dtp & DTR  |  dtn & dtp & dtr  ; 
assign FGF = ~fgf;  //complement 
assign FFA =  DTA & dtc & dte  |  dta & DTC & dte  |  dta & dtc & DTE  |  DTA & DTC & DTE  ; 
assign ffa = ~FFA; //complement 
assign ffb =  DTA & dtc & dte  |  dta & DTC & dte  |  dta & dtc & DTE  |  dta & dtc & dte  ; 
assign FFB = ~ffb;  //complement 
assign dgj = ~DGJ;  //complement 
assign DGK = ~dgk;  //complement 
assign abl = ~ABL;  //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign FFC =  DTG & dti & dtk  |  dtg & DTI & dtk  |  dtg & dti & DTK  |  DTG & DTI & DTK  ; 
assign ffc = ~FFC; //complement 
assign ffd =  DTG & dti & dtk  |  dtg & DTI & dtk  |  dtg & dti & DTK  |  dtg & dti & dtk  ; 
assign FFD = ~ffd;  //complement 
assign FFE =  DTM & dto & dtq  |  dtm & DTO & dtq  |  dtm & dto & DTQ  |  DTM & DTO & DTQ  ; 
assign ffe = ~FFE; //complement 
assign fff =  DTM & dto & dtq  |  dtm & DTO & dtq  |  dtm & dto & DTQ  |  dtm & dto & dtq  ; 
assign FFF = ~fff;  //complement 
assign dha = ~DHA;  //complement 
assign DHB = ~dhb;  //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign FEA =  DSB & dsd & dsf  |  dsb & DSD & dsf  |  dsb & dsd & DSF  |  DSB & DSD & DSF  ; 
assign fea = ~FEA; //complement 
assign feb =  DSB & dsd & dsf  |  dsb & DSD & dsf  |  dsb & dsd & DSF  |  dsb & dsd & dsf  ; 
assign FEB = ~feb;  //complement 
assign FEC =  DSH & dsj & dsl  |  dsh & DSJ & dsl  |  dsh & dsj & DSL  |  DSH & DSJ & DSL  ; 
assign fec = ~FEC; //complement 
assign fed =  DSH & dsj & dsl  |  dsh & DSJ & dsl  |  dsh & dsj & DSL  |  dsh & dsj & dsl  ; 
assign FED = ~fed;  //complement 
assign dhc = ~DHC;  //complement 
assign DHD = ~dhd;  //complement 
assign gld = ~GLD;  //complement 
assign FEE =  DSN & dsp & dsr  |  dsn & DSP & dsr  |  dsn & dsp & DSR  |  DSN & DSP & DSR  ; 
assign fee = ~FEE; //complement 
assign fef =  DSN & dsp & dsr  |  dsn & DSP & dsr  |  dsn & dsp & DSR  |  dsn & dsp & dsr  ; 
assign FEF = ~fef;  //complement 
assign FDA =  DSA & dsc & dse  |  dsa & DSC & dse  |  dsa & dsc & DSE  |  DSA & DSC & DSE  ; 
assign fda = ~FDA; //complement 
assign fdb =  DSA & dsc & dse  |  dsa & DSC & dse  |  dsa & dsc & DSE  |  dsa & dsc & dse  ; 
assign FDB = ~fdb;  //complement 
assign dia = ~DIA;  //complement 
assign DIB = ~dib;  //complement 
assign drs = ~DRS;  //complement 
assign gbe = ~GBE;  //complement 
assign gce = ~GCE;  //complement 
assign gde = ~GDE;  //complement 
assign FDC =  DSG & dsi & dsk  |  dsg & DSI & dsk  |  dsg & dsi & DSK  |  DSG & DSI & DSK  ; 
assign fdc = ~FDC; //complement 
assign fdd =  DSG & dsi & dsk  |  dsg & DSI & dsk  |  dsg & dsi & DSK  |  dsg & dsi & dsk  ; 
assign FDD = ~fdd;  //complement 
assign FDE =  DSM & dso & dsq  |  dsm & DSO & dsq  |  dsm & dso & DSQ  |  DSM & DSO & DSQ  ; 
assign fde = ~FDE; //complement 
assign fdf =  DSM & dso & dsq  |  dsm & DSO & dsq  |  dsm & dso & DSQ  |  dsm & dso & dsq  ; 
assign FDF = ~fdf;  //complement 
assign dic = ~DIC;  //complement 
assign DID = ~did;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign abc = ~ABC;  //complement 
assign FCA =  DRB & drd & drf  |  drb & DRD & drf  |  drb & drd & DRF  |  DRB & DRD & DRF  ; 
assign fca = ~FCA; //complement 
assign fcb =  DRB & drd & drf  |  drb & DRD & drf  |  drb & drd & DRF  |  drb & drd & drf  ; 
assign FCB = ~fcb;  //complement 
assign FCC =  DRH & drj & drl  |  drh & DRJ & drl  |  drh & drj & DRL  |  DRH & DRJ & DRL  ; 
assign fcc = ~FCC; //complement 
assign fcd =  DRH & drj & drl  |  drh & DRJ & drl  |  drh & drj & DRL  |  drh & drj & drl  ; 
assign FCD = ~fcd;  //complement 
assign die = ~DIE;  //complement 
assign DIF = ~dif;  //complement 
assign abd = ~ABD;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign FCE =  DRN & drp & drr  |  drn & DRP & drr  |  drn & drp & DRR  |  DRN & DRP & DRR  ; 
assign fce = ~FCE; //complement 
assign fcf =  DRN & drp & drr  |  drn & DRP & drr  |  drn & drp & DRR  |  drn & drp & drr  ; 
assign FCF = ~fcf;  //complement 
assign FBA =  DRA & drc & dre  |  dra & DRC & dre  |  dra & drc & DRE  |  DRA & DRC & DRE  ; 
assign fba = ~FBA; //complement 
assign fbb =  DRA & drc & dre  |  dra & DRC & dre  |  dra & drc & DRE  |  dra & drc & dre  ; 
assign FBB = ~fbb;  //complement 
assign CAA =  BAA & ACA  ; 
assign caa = ~CAA;  //complement 
assign CAB =  BAA & ACC  ; 
assign cab = ~CAB;  //complement 
assign CAC =  BAA & ACE  ; 
assign cac = ~CAC;  //complement 
assign CPB =  BAP & ACB  ; 
assign cpb = ~CPB;  //complement 
assign CPC =  BAP & ACD  ; 
assign cpc = ~CPC;  //complement 
assign CPD =  BAP & ACF  ; 
assign cpd = ~CPD;  //complement 
assign baa = ~BAA;  //complement 
assign bab = ~BAB;  //complement 
assign bac = ~BAC;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign oac = ~OAC;  //complement 
assign CAD =  BAA & ACG  ; 
assign cad = ~CAD;  //complement 
assign CAE =  BAA & ACI  ; 
assign cae = ~CAE;  //complement 
assign CAF =  BAA & ACK  ; 
assign caf = ~CAF;  //complement 
assign CPE =  BAP & ACH  ; 
assign cpe = ~CPE;  //complement 
assign CPF =  BAP & ACJ  ; 
assign cpf = ~CPF;  //complement 
assign CPG =  BAP & ACL  ; 
assign cpg = ~CPG;  //complement 
assign bad = ~BAD;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign oad = ~OAD;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign CAG =  BAA & ACM  ; 
assign cag = ~CAG;  //complement 
assign CAH =  BAA & ACO  ; 
assign cah = ~CAH;  //complement 
assign CAI =  BAA & ADA  ; 
assign cai = ~CAI;  //complement 
assign CPH =  BAP & ACN  ; 
assign cph = ~CPH;  //complement 
assign CPI =  BAP & ACP  ; 
assign cpi = ~CPI;  //complement 
assign CQA =  BBA & ACA  ; 
assign cqa = ~CQA;  //complement 
assign bai = ~BAI;  //complement 
assign baj = ~BAJ;  //complement 
assign bak = ~BAK;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign CAJ =  BAA & ADC  ; 
assign caj = ~CAJ;  //complement 
assign CAK =  BAA & ADE  ; 
assign cak = ~CAK;  //complement 
assign CAL =  BAA & ADG  ; 
assign cal = ~CAL;  //complement 
assign CQB =  BBA & ACC  ; 
assign cqb = ~CQB;  //complement 
assign CQC =  BBA & ACE  ; 
assign cqc = ~CQC;  //complement 
assign CQD =  BBA & ACG  ; 
assign cqd = ~CQD;  //complement 
assign bal = ~BAL;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign oak = ~OAK;  //complement 
assign CAM =  BAA & ADI  ; 
assign cam = ~CAM;  //complement 
assign CAN =  BAA & ADK  ; 
assign can = ~CAN;  //complement 
assign CAO =  BAA & ADM  ; 
assign cao = ~CAO;  //complement 
assign CQE =  BBA & ACI  ; 
assign cqe = ~CQE;  //complement 
assign CQF =  BBA & ACK  ; 
assign cqf = ~CQF;  //complement 
assign CQG =  BBA & ACM  ; 
assign cqg = ~CQG;  //complement 
assign bbi = ~BBI;  //complement 
assign bbj = ~BBJ;  //complement 
assign bbk = ~BBK;  //complement 
assign oal = ~OAL;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign CAP =  BAA & ADO  ; 
assign cap = ~CAP;  //complement 
assign CBA =  BAB & ACQ  ; 
assign cba = ~CBA;  //complement 
assign CBB =  BAB & ACB  ; 
assign cbb = ~CBB;  //complement 
assign CQH =  BBA & ACO  ; 
assign cqh = ~CQH;  //complement 
assign CRA =  BBB & ACQ  ; 
assign cra = ~CRA;  //complement 
assign CRB =  BBB & ACB  ; 
assign crb = ~CRB;  //complement 
assign bbl = ~BBL;  //complement 
assign bbm = ~BBM;  //complement 
assign bbn = ~BBN;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign CBC =  BAB & ACD  ; 
assign cbc = ~CBC;  //complement 
assign CBD =  BAB & ACF  ; 
assign cbd = ~CBD;  //complement 
assign CBE =  BAB & ACH  ; 
assign cbe = ~CBE;  //complement 
assign CRC =  BBB & ACD  ; 
assign crc = ~CRC;  //complement 
assign CRD =  BBB & ACF  ; 
assign crd = ~CRD;  //complement 
assign CRE =  BBB & ACH  ; 
assign cre = ~CRE;  //complement 
assign dgf = ~DGF;  //complement 
assign dlk = ~DLK;  //complement 
assign doo = ~DOO;  //complement 
assign pal = ~PAL;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign obc = ~OBC;  //complement 
assign CBF =  BAB & ACJ  ; 
assign cbf = ~CBF;  //complement 
assign CBG =  BAB & ACL  ; 
assign cbg = ~CBG;  //complement 
assign CBH =  BAB & ACN  ; 
assign cbh = ~CBH;  //complement 
assign CRF =  BBB & ACJ  ; 
assign crf = ~CRF;  //complement 
assign CRG =  BBB & ACL  ; 
assign crg = ~CRG;  //complement 
assign CRH =  BBB & ACN  ; 
assign crh = ~CRH;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign obg = ~OBG;  //complement 
assign obd = ~OBD;  //complement 
assign EPD =  DLH & DLJ  ; 
assign epd = ~EPD;  //complement 
assign NKB =  NFA  ; 
assign nkb = ~NKB;  //complement 
assign END =  DKH & DKJ  ; 
assign end = ~END;  //complement 
assign NEE = ~nee;  //complement 
assign mbf = ~MBF;  //complement 
assign MDF = ~mdf;  //complement 
assign dso = ~DSO;  //complement 
assign DSP = ~dsp;  //complement 
assign NEF = ~nef;  //complement 
assign NEG = ~neg;  //complement 
assign mbg = ~MBG;  //complement 
assign MDG = ~mdg;  //complement 
assign dsq = ~DSQ;  //complement 
assign DSR = ~dsr;  //complement 
assign dhe = ~DHE;  //complement 
assign neh = ~NEH;  //complement 
assign mbh = ~MBH;  //complement 
assign MDH = ~mdh;  //complement 
assign dss = ~DSS;  //complement 
assign DST = ~dst;  //complement 
assign NEI = ~nei;  //complement 
assign NEJ = ~nej;  //complement 
assign NEK = ~nek;  //complement 
assign dta = ~DTA;  //complement 
assign DTB = ~dtb;  //complement 
assign dtu = ~DTU;  //complement 
assign dtv = ~DTV;  //complement 
assign FFG =  DTS & dtu  |  dts & DTU  ; 
assign ffg = ~FFG;  //complement 
assign dtc = ~DTC;  //complement 
assign DTD = ~dtd;  //complement 
assign FGG =  DTT & dtv  |  dtt & DTV  ; 
assign fgg = ~FGG;  //complement 
assign EUF =  DOM & DOO  ; 
assign euf = ~EUF;  //complement 
assign EXF =  DPN & DPP  ; 
assign exf = ~EXF;  //complement 
assign FGH =  DTT & DTV  ; 
assign fgh = ~FGH;  //complement 
assign EWF = DPO & DPM ; 
assign ewf = ~EWF ; //complement 
assign dte = ~DTE;  //complement 
assign DTF = ~dtf;  //complement 
assign EIC = DIG; 
assign eic = ~EIC; //complement 
assign HGC = GHD; 
assign hgc = ~HGC;  //complement 
assign nub = nbi; 
assign NUB = ~nub;  //complement 
assign nvb = nbm; 
assign NVB = ~nvb;  //complement 
assign ECA =  DGD & dgf  |  dgd & DGF  ; 
assign eca = ~ECA;  //complement 
assign EEA =  DGG & dgj  |  dgg & DGJ  ; 
assign eea = ~EEA;  //complement 
assign EMC =  DKG & dki  |  dkg & DKI  ; 
assign emc = ~EMC;  //complement 
assign EPC =  DLH & dlj  |  dlh & DLJ  ; 
assign epc = ~EPC;  //complement 
assign EXE =  DPN & dpp  |  dpn & DPP  ; 
assign exe = ~EXE;  //complement 
assign bbd = ~BBD;  //complement 
assign bbe = ~BBE;  //complement 
assign bbf = ~BBF;  //complement 
assign bba = ~BBA;  //complement 
assign bbb = ~BBB;  //complement 
assign bbc = ~BBC;  //complement 
assign dtg = ~DTG;  //complement 
assign DTH = ~dth;  //complement 
assign dti = ~DTI;  //complement 
assign DTJ = ~dtj;  //complement 
assign dja = ~DJA;  //complement 
assign DJB = ~djb;  //complement 
assign gzm = ~GZM;  //complement 
assign FBC =  DRG & dri & drk  |  drg & DRI & drk  |  drg & dri & DRK  |  DRG & DRI & DRK  ; 
assign fbc = ~FBC; //complement 
assign fbd =  DRG & dri & drk  |  drg & DRI & drk  |  drg & dri & DRK  |  drg & dri & drk  ; 
assign FBD = ~fbd;  //complement 
assign FBE =  DRM & dro & drq  |  drm & DRO & drq  |  drm & dro & DRQ  |  DRM & DRO & DRQ  ; 
assign fbe = ~FBE; //complement 
assign fbf =  DRM & dro & drq  |  drm & DRO & drq  |  drm & dro & DRQ  |  drm & dro & drq  ; 
assign FBF = ~fbf;  //complement 
assign djc = ~DJC;  //complement 
assign DJD = ~djd;  //complement 
assign NEL = ~nel;  //complement 
assign FAA =  DQB & dqd & dqf  |  dqb & DQD & dqf  |  dqb & dqd & DQF  |  DQB & DQD & DQF  ; 
assign faa = ~FAA; //complement 
assign fab =  DQB & dqd & dqf  |  dqb & DQD & dqf  |  dqb & dqd & DQF  |  dqb & dqd & dqf  ; 
assign FAB = ~fab;  //complement 
assign FAC =  DQH & dqj & dql  |  dqh & DQJ & dql  |  dqh & dqj & DQL  |  DQH & DQJ & DQL  ; 
assign fac = ~FAC; //complement 
assign fad =  DQH & dqj & dql  |  dqh & DQJ & dql  |  dqh & dqj & DQL  |  dqh & dqj & dql  ; 
assign FAD = ~fad;  //complement 
assign dje = ~DJE;  //complement 
assign DJF = ~djf;  //complement 
assign NEM = ~nem;  //complement 
assign FAE =  DQN & dqp & dqr  |  dqn & DQP & dqr  |  dqn & dqp & DQR  |  DQN & DQP & DQR  ; 
assign fae = ~FAE; //complement 
assign faf =  DQN & dqp & dqr  |  dqn & DQP & dqr  |  dqn & dqp & DQR  |  dqn & dqp & dqr  ; 
assign FAF = ~faf;  //complement 
assign EYA =  DQA & dqc & dqe  |  dqa & DQC & dqe  |  dqa & dqc & DQE  |  DQA & DQC & DQE  ; 
assign eya = ~EYA; //complement 
assign eyb =  DQA & dqc & dqe  |  dqa & DQC & dqe  |  dqa & dqc & DQE  |  dqa & dqc & dqe  ; 
assign EYB = ~eyb;  //complement 
assign djg = ~DJG;  //complement 
assign DJH = ~djh;  //complement 
assign HAC =  GBB & gbd  |  gbb & GBD  ; 
assign hac = ~HAC;  //complement 
assign EYC =  DQG & dqi & dqk  |  dqg & DQI & dqk  |  dqg & dqi & DQK  |  DQG & DQI & DQK  ; 
assign eyc = ~EYC; //complement 
assign eyd =  DQG & dqi & dqk  |  dqg & DQI & dqk  |  dqg & dqi & DQK  |  dqg & dqi & dqk  ; 
assign EYD = ~eyd;  //complement 
assign EYE =  DQM & dqo & dqq  |  dqm & DQO & dqq  |  dqm & dqo & DQQ  |  DQM & DQO & DQQ  ; 
assign eye = ~EYE; //complement 
assign eyf =  DQM & dqo & dqq  |  dqm & DQO & dqq  |  dqm & dqo & DQQ  |  dqm & dqo & dqq  ; 
assign EYF = ~eyf;  //complement 
assign dka = ~DKA;  //complement 
assign DKB = ~dkb;  //complement 
assign HBC =  GCB & gcd  |  gcb & GCD  ; 
assign hbc = ~HBC;  //complement 
assign EXA =  DPB & dpd & dpf  |  dpb & DPD & dpf  |  dpb & dpd & DPF  |  DPB & DPD & DPF  ; 
assign exa = ~EXA; //complement 
assign exb =  DPB & dpd & dpf  |  dpb & DPD & dpf  |  dpb & dpd & DPF  |  dpb & dpd & dpf  ; 
assign EXB = ~exb;  //complement 
assign EXC =  DPH & dpj & dpl  |  dph & DPJ & dpl  |  dph & dpj & DPL  |  DPH & DPJ & DPL  ; 
assign exc = ~EXC; //complement 
assign exd =  DPH & dpj & dpl  |  dph & DPJ & dpl  |  dph & dpj & DPL  |  dph & dpj & dpl  ; 
assign EXD = ~exd;  //complement 
assign dkc = ~DKC;  //complement 
assign DKD = ~dkd;  //complement 
assign HCD =  GDB & gdd  |  gdb & GDD  ; 
assign hcd = ~HCD;  //complement 
assign EWA =  DPA & dpc & dpe  |  dpa & DPC & dpe  |  dpa & dpc & DPE  |  DPA & DPC & DPE  ; 
assign ewa = ~EWA; //complement 
assign ewb =  DPA & dpc & dpe  |  dpa & DPC & dpe  |  dpa & dpc & DPE  |  dpa & dpc & dpe  ; 
assign EWB = ~ewb;  //complement 
assign EWC =  DPG & dpi & dpk  |  dpg & DPI & dpk  |  dpg & dpi & DPK  |  DPG & DPI & DPK  ; 
assign ewc = ~EWC; //complement 
assign ewd =  DPG & dpi & dpk  |  dpg & DPI & dpk  |  dpg & dpi & DPK  |  dpg & dpi & dpk  ; 
assign EWD = ~ewd;  //complement 
assign dke = ~DKE;  //complement 
assign DKF = ~dkf;  //complement 
assign gnd = ~GND;  //complement 
assign EWE =  DPM & dpo  |  dpm & DPO  ; 
assign ewe = ~EWE;  //complement 
assign EVA =  DOB & dod & dof  |  dob & DOD & dof  |  dob & dod & DOF  |  DOB & DOD & DOF  ; 
assign eva = ~EVA; //complement 
assign evb =  DOB & dod & dof  |  dob & DOD & dof  |  dob & dod & DOF  |  dob & dod & dof  ; 
assign EVB = ~evb;  //complement 
assign dkg = ~DKG;  //complement 
assign DKH = ~dkh;  //complement 
assign gzf = ~GZF;  //complement 
assign EVC =  DOH & doj & dol  |  doh & DOJ & dol  |  doh & doj & DOL  |  DOH & DOJ & DOL  ; 
assign evc = ~EVC; //complement 
assign evd =  DOH & doj & dol  |  doh & DOJ & dol  |  doh & doj & DOL  |  doh & doj & dol  ; 
assign EVD = ~evd;  //complement 
assign EUA =  DOA & doc & doe  |  doa & DOC & doe  |  doa & doc & DOE  |  DOA & DOC & DOE  ; 
assign eua = ~EUA; //complement 
assign eub =  DOA & doc & doe  |  doa & DOC & doe  |  doa & doc & DOE  |  doa & doc & doe  ; 
assign EUB = ~eub;  //complement 
assign CBI =  BAB & ACP  ; 
assign cbi = ~CBI;  //complement 
assign CBJ =  BAB & ADB  ; 
assign cbj = ~CBJ;  //complement 
assign CBK =  BAB & ADD  ; 
assign cbk = ~CBK;  //complement 
assign CSA =  BBC & ACA  ; 
assign csa = ~CSA;  //complement 
assign CSB =  BBC & ACC  ; 
assign csb = ~CSB;  //complement 
assign CSC =  BBC & ACE  ; 
assign csc = ~CSC;  //complement 
assign gfe = ~GFE;  //complement 
assign ghe = ~GHE;  //complement 
assign goc = ~GOC;  //complement 
assign gpc = ~GPC;  //complement 
assign obh = ~OBH;  //complement 
assign CBL =  BAB & ADF  ; 
assign cbl = ~CBL;  //complement 
assign CBM =  BAB & ADH  ; 
assign cbm = ~CBM;  //complement 
assign CBN =  BAB & ADJ  ; 
assign cbn = ~CBN;  //complement 
assign CSD =  BBC & ACG  ; 
assign csd = ~CSD;  //complement 
assign CSE =  BBC & ACI  ; 
assign cse = ~CSE;  //complement 
assign CSF =  BBC & ACK  ; 
assign csf = ~CSF;  //complement 
assign gqc = ~GQC;  //complement 
assign gzk = ~GZK;  //complement 
assign gzl = ~GZL;  //complement 
assign gzh = ~GZH;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign obk = ~OBK;  //complement 
assign CBO =  BAB & ADL  ; 
assign cbo = ~CBO;  //complement 
assign CBP =  BAB & ADN  ; 
assign cbp = ~CBP;  //complement 
assign CCA =  BAC & ACA  ; 
assign cca = ~CCA;  //complement 
assign CSG =  BBC & ACM  ; 
assign csg = ~CSG;  //complement 
assign CTA =  BBD & ACQ  ; 
assign cta = ~CTA;  //complement 
assign CTB =  BBD & ACB  ; 
assign ctb = ~CTB;  //complement 
assign HZG = GZM; 
assign hzg = ~HZG; //complement 
assign HZI = GZH; 
assign hzi = ~HZI;  //complement 
assign HZK = GZK; 
assign hzk = ~HZK;  //complement 
assign obl = ~OBL;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign CCB =  BAC & ACC  ; 
assign ccb = ~CCB;  //complement 
assign CCC =  BAC & ACE  ; 
assign ccc = ~CCC;  //complement 
assign CCD =  BAC & ACG  ; 
assign ccd = ~CCD;  //complement 
assign CTC =  BBD & ACD  ; 
assign ctc = ~CTC;  //complement 
assign CTD =  BBD & ACF  ; 
assign ctd = ~CTD;  //complement 
assign CTE =  BBD & ACH  ; 
assign cte = ~CTE;  //complement 
assign jac = ~JAC;  //complement 
assign jbc = ~JBC;  //complement 
assign jcc = ~JCC;  //complement 
assign dig = ~DIG;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign CCE =  BAC & ACI  ; 
assign cce = ~CCE;  //complement 
assign CCF =  BAC & ACK  ; 
assign ccf = ~CCF;  //complement 
assign CCG =  BAC & ACM  ; 
assign ccg = ~CCG;  //complement 
assign CTF =  BBD & ACJ  ; 
assign ctf = ~CTF;  //complement 
assign CTG =  BBD & ACL  ; 
assign ctg = ~CTG;  //complement 
assign CUA =  BBE & ACA  ; 
assign cua = ~CUA;  //complement 
assign jec = ~JEC;  //complement 
assign jgc = ~JGC;  //complement 
assign HBD =  GCB & GCD  ; 
assign hbd = ~HBD;  //complement 
assign HZF =  GZF & GZN  ; 
assign hzf = ~HZF;  //complement 
assign HCE =  GDB & GDD  ; 
assign hce = ~HCE;  //complement 
assign CCH =  BAC & ACO  ; 
assign cch = ~CCH;  //complement 
assign CCI =  BAC & ADA  ; 
assign cci = ~CCI;  //complement 
assign CCJ =  BAC & ADC  ; 
assign ccj = ~CCJ;  //complement 
assign CUB =  BBE & ACC  ; 
assign cub = ~CUB;  //complement 
assign CUC =  BBE & ACE  ; 
assign cuc = ~CUC;  //complement 
assign CUD =  BBE & ACG  ; 
assign cud = ~CUD;  //complement 
assign jzg = ~JZG;  //complement 
assign jzi = ~JZI;  //complement 
assign jzk = ~JZK;  //complement 
assign jzl = ~JZL;  //complement 
assign NEO = ~neo;  //complement 
assign CCK =  BAC & ADE  ; 
assign cck = ~CCK;  //complement 
assign CCL =  BAC & ADG  ; 
assign ccl = ~CCL;  //complement 
assign CCM =  BAC & ADI  ; 
assign ccm = ~CCM;  //complement 
assign CUE =  BBE & ACI  ; 
assign cue = ~CUE;  //complement 
assign CUF =  BBE & ACK  ; 
assign cuf = ~CUF;  //complement 
assign CVA =  BBF & ACQ  ; 
assign cva = ~CVA;  //complement 
assign gmd = ~GMD;  //complement 
assign kba = ~KBA;  //complement 
assign KBB = ~kbb;  //complement 
assign kbc = ~KBC;  //complement 
assign kca = ~KCA;  //complement 
assign CCN =  BAC & ADK  ; 
assign ccn = ~CCN;  //complement 
assign CCO =  BAC & ADM  ; 
assign cco = ~CCO;  //complement 
assign CDA =  BAD & ACQ  ; 
assign cda = ~CDA;  //complement 
assign CVB =  BBF & ACB  ; 
assign cvb = ~CVB;  //complement 
assign CVC =  BBF & ACD  ; 
assign cvc = ~CVC;  //complement 
assign CVD =  BBF & ACF  ; 
assign cvd = ~CVD;  //complement 
assign KCB = ~kcb;  //complement 
assign kcc = ~KCC;  //complement 
assign kda = ~KDA;  //complement 
assign KDB = ~kdb;  //complement 
assign NEN = ~nen;  //complement 
assign aaq = ~AAQ;  //complement 
assign gfc = ~GFC;  //complement 
assign GFD = ~gfd;  //complement 
assign gbc = ~GBC;  //complement 
assign GBD = ~gbd;  //complement 
assign dtk = ~DTK;  //complement 
assign DTL = ~dtl;  //complement 
assign NEP = ~nep;  //complement 
assign gga = ~GGA;  //complement 
assign GGB = ~ggb;  //complement 
assign gca = ~GCA;  //complement 
assign GCB = ~gcb;  //complement 
assign dtm = ~DTM;  //complement 
assign DTN = ~dtn;  //complement 
assign gzd = ~GZD;  //complement 
assign ggc = ~GGC;  //complement 
assign GGD = ~ggd;  //complement 
assign gcc = ~GCC;  //complement 
assign GCD = ~gcd;  //complement 
assign dto = ~DTO;  //complement 
assign DTP = ~dtp;  //complement 
assign dhf = ~DHF;  //complement 
assign gha = ~GHA;  //complement 
assign GHB = ~ghb;  //complement 
assign gda = ~GDA;  //complement 
assign GDB = ~gdb;  //complement 
assign dtq = ~DTQ;  //complement 
assign DTR = ~dtr;  //complement 
assign LFC =  KGB & kfc  |  kgb & KFC  ; 
assign lfc = ~LFC;  //complement 
assign ghc = ~GHC;  //complement 
assign GHD = ~ghd;  //complement 
assign gdc = ~GDC;  //complement 
assign GDD = ~gdd;  //complement 
assign dts = ~DTS;  //complement 
assign DTT = ~dtt;  //complement 
assign gmc = ~GMC;  //complement 
assign gia = ~GIA;  //complement 
assign GIB = ~gib;  //complement 
assign gea = ~GEA;  //complement 
assign GEB = ~geb;  //complement 
assign gaa = ~GAA;  //complement 
assign GAB = ~gab;  //complement 
assign HDC =  GEB & ged  |  geb & GED  ; 
assign hdc = ~HDC;  //complement 
assign gec = ~GEC;  //complement 
assign GED = ~ged;  //complement 
assign HDD = GED & GEB ; 
assign hdd = ~HDD ; //complement 
assign gfa = ~GFA;  //complement 
assign GFB = ~gfb;  //complement 
assign gic = ~GIC;  //complement 
assign GID = ~gid;  //complement 
assign gja = ~GJA;  //complement 
assign GJB = ~gjb;  //complement 
assign gac = ~GAC;  //complement 
assign GAD = ~gad;  //complement 
assign gba = ~GBA;  //complement 
assign GBB = ~gbb;  //complement 
assign dla = ~DLA;  //complement 
assign DLB = ~dlb;  //complement 
assign OIA = ~oia;  //complement 
assign OKA = ~oka;  //complement 
assign OMA = ~oma;  //complement 
assign OOA = ~ooa;  //complement 
assign EUC =  DOG & doi & dok  |  dog & DOI & dok  |  dog & doi & DOK  |  DOG & DOI & DOK  ; 
assign euc = ~EUC; //complement 
assign eud =  DOG & doi & dok  |  dog & DOI & dok  |  dog & doi & DOK  |  dog & doi & dok  ; 
assign EUD = ~eud;  //complement 
assign ETA =  DNB & dnd & dnf  |  dnb & DND & dnf  |  dnb & dnd & DNF  |  DNB & DND & DNF  ; 
assign eta = ~ETA; //complement 
assign etb =  DNB & dnd & dnf  |  dnb & DND & dnf  |  dnb & dnd & DNF  |  dnb & dnd & dnf  ; 
assign ETB = ~etb;  //complement 
assign dlc = ~DLC;  //complement 
assign DLD = ~dld;  //complement 
assign NFA = ~nfa;  //complement 
assign ETC =  DNH & dnj & dnl  |  dnh & DNJ & dnl  |  dnh & dnj & DNL  |  DNH & DNJ & DNL  ; 
assign etc = ~ETC; //complement 
assign etd =  DNH & dnj & dnl  |  dnh & DNJ & dnl  |  dnh & dnj & DNL  |  dnh & dnj & dnl  ; 
assign ETD = ~etd;  //complement 
assign ESA =  DNA & dnc & dne  |  dna & DNC & dne  |  dna & dnc & DNE  |  DNA & DNC & DNE  ; 
assign esa = ~ESA; //complement 
assign esb =  DNA & dnc & dne  |  dna & DNC & dne  |  dna & dnc & DNE  |  dna & dnc & dne  ; 
assign ESB = ~esb;  //complement 
assign dle = ~DLE;  //complement 
assign DLF = ~dlf;  //complement 
assign NTD =  NBE & NBF & NBG  |  NBG & NFF  |  NFG  ; 
assign ntd = ~NTD; //complement 
assign ESC =  DNG & dni & dnk  |  dng & DNI & dnk  |  dng & dni & DNK  |  DNG & DNI & DNK  ; 
assign esc = ~ESC; //complement 
assign esd =  DNG & dni & dnk  |  dng & DNI & dnk  |  dng & dni & DNK  |  dng & dni & dnk  ; 
assign ESD = ~esd;  //complement 
assign ERA =  DMB & dmd & dmf  |  dmb & DMD & dmf  |  dmb & dmd & DMF  |  DMB & DMD & DMF  ; 
assign era = ~ERA; //complement 
assign erb =  DMB & dmd & dmf  |  dmb & DMD & dmf  |  dmb & dmd & DMF  |  dmb & dmd & dmf  ; 
assign ERB = ~erb;  //complement 
assign dlg = ~DLG;  //complement 
assign DLH = ~dlh;  //complement 
assign glc = ~GLC;  //complement 
assign ERC =  DMH & dmj & dml  |  dmh & DMJ & dml  |  dmh & dmj & DML  |  DMH & DMJ & DML  ; 
assign erc = ~ERC; //complement 
assign erd =  DMH & dmj & dml  |  dmh & DMJ & dml  |  dmh & dmj & DML  |  dmh & dmj & dml  ; 
assign ERD = ~erd;  //complement 
assign EQA =  DMA & dmc & dme  |  dma & DMC & dme  |  dma & dmc & DME  |  DMA & DMC & DME  ; 
assign eqa = ~EQA; //complement 
assign eqb =  DMA & dmc & dme  |  dma & DMC & dme  |  dma & dmc & DME  |  dma & dmc & dme  ; 
assign EQB = ~eqb;  //complement 
assign dli = ~DLI;  //complement 
assign DLJ = ~dlj;  //complement 
assign HAD =  GBB & GBD  ; 
assign had = ~HAD;  //complement 
assign nrb =  nam  ; 
assign NRB = ~nrb;  //complement 
assign FDG =  DSS  ; 
assign fdg = ~FDG;  //complement 
assign EQC =  DMG & dmi & dmk  |  dmg & DMI & dmk  |  dmg & dmi & DMK  |  DMG & DMI & DMK  ; 
assign eqc = ~EQC; //complement 
assign eqd =  DMG & dmi & dmk  |  dmg & DMI & dmk  |  dmg & dmi & DMK  |  dmg & dmi & dmk  ; 
assign EQD = ~eqd;  //complement 
assign EPA =  DLB & dld & dlf  |  dlb & DLD & dlf  |  dlb & dld & DLF  |  DLB & DLD & DLF  ; 
assign epa = ~EPA; //complement 
assign epb =  DLB & dld & dlf  |  dlb & DLD & dlf  |  dlb & dld & DLF  |  dlb & dld & dlf  ; 
assign EPB = ~epb;  //complement 
assign dma = ~DMA;  //complement 
assign DMB = ~dmb;  //complement 
assign mbj = ~MBJ;  //complement 
assign EOA =  DLA & dlc & dle  |  dla & DLC & dle  |  dla & dlc & DLE  |  DLA & DLC & DLE  ; 
assign eoa = ~EOA; //complement 
assign eob =  DLA & dlc & dle  |  dla & DLC & dle  |  dla & dlc & DLE  |  dla & dlc & dle  ; 
assign EOB = ~eob;  //complement 
assign EOC =  DLG & dli & dlk  |  dlg & DLI & dlk  |  dlg & dli & DLK  |  DLG & DLI & DLK  ; 
assign eoc = ~EOC; //complement 
assign eod =  DLG & dli & dlk  |  dlg & DLI & dlk  |  dlg & dli & DLK  |  dlg & dli & dlk  ; 
assign EOD = ~eod;  //complement 
assign dmc = ~DMC;  //complement 
assign DMD = ~dmd;  //complement 
assign mec = ~MEC;  //complement 
assign ENA =  DKB & dkd & dkf  |  dkb & DKD & dkf  |  dkb & dkd & DKF  |  DKB & DKD & DKF  ; 
assign ena = ~ENA; //complement 
assign enb =  DKB & dkd & dkf  |  dkb & DKD & dkf  |  dkb & dkd & DKF  |  dkb & dkd & dkf  ; 
assign ENB = ~enb;  //complement 
assign EMA =  DKA & dkc & dke  |  dka & DKC & dke  |  dka & dkc & DKE  |  DKA & DKC & DKE  ; 
assign ema = ~EMA; //complement 
assign emb =  DKA & dkc & dke  |  dka & DKC & dke  |  dka & dkc & DKE  |  dka & dkc & dke  ; 
assign EMB = ~emb;  //complement 
assign dme = ~DME;  //complement 
assign DMF = ~dmf;  //complement 
assign OIH = ~oih;  //complement 
assign OKH = ~okh;  //complement 
assign OMH = ~omh;  //complement 
assign OOH = ~ooh;  //complement 
assign ELA =  DJB & djd & djf  |  djb & DJD & djf  |  djb & djd & DJF  |  DJB & DJD & DJF  ; 
assign ela = ~ELA; //complement 
assign elb =  DJB & djd & djf  |  djb & DJD & djf  |  djb & djd & DJF  |  djb & djd & djf  ; 
assign ELB = ~elb;  //complement 
assign EKA =  DJA & dje & djc  |  dja & DJE & djc  |  dja & dje & DJC  |  DJA & DJE & DJC  ; 
assign eka = ~EKA; //complement 
assign ekb =  DJA & dje & djc  |  dja & DJE & djc  |  dja & dje & DJC  |  dja & dje & djc  ; 
assign EKB = ~ekb;  //complement 
assign CDB =  BAD & ACB  ; 
assign cdb = ~CDB;  //complement 
assign CDC =  BAD & ACD  ; 
assign cdc = ~CDC;  //complement 
assign CDD =  BAD & ACF  ; 
assign cdd = ~CDD;  //complement 
assign CVE =  BBF & ACH  ; 
assign cve = ~CVE;  //complement 
assign CVF =  BBF & ACJ  ; 
assign cvf = ~CVF;  //complement 
assign CWA =  BBG & ACA  ; 
assign cwa = ~CWA;  //complement 
assign kdc = ~KDC;  //complement 
assign kea = ~KEA;  //complement 
assign KEB = ~keb;  //complement 
assign kfc = ~KFC;  //complement 
assign gjc = ~GJC;  //complement 
assign CDE =  BAD & ACH  ; 
assign cde = ~CDE;  //complement 
assign CDF =  BAD & ACJ  ; 
assign cdf = ~CDF;  //complement 
assign CDG =  BAD & ACL  ; 
assign cdg = ~CDG;  //complement 
assign CWB =  BBG & ACC  ; 
assign cwb = ~CWB;  //complement 
assign CWC =  BBG & ACE  ; 
assign cwc = ~CWC;  //complement 
assign CWD =  BBG & ACG  ; 
assign cwd = ~CWD;  //complement 
assign kfa = ~KFA;  //complement 
assign KFB = ~kfb;  //complement 
assign kga = ~KGA;  //complement 
assign KGB = ~kgb;  //complement 
assign mbk = ~MBK;  //complement 
assign CDH =  BAD & ACN  ; 
assign cdh = ~CDH;  //complement 
assign CDI =  BAD & ACP  ; 
assign cdi = ~CDI;  //complement 
assign CDJ =  BAD & ADB  ; 
assign cdj = ~CDJ;  //complement 
assign CWE =  BBG & ACI  ; 
assign cwe = ~CWE;  //complement 
assign CXA =  BBH & ACQ  ; 
assign cxa = ~CXA;  //complement 
assign CXB =  BBH & ACB  ; 
assign cxb = ~CXB;  //complement 
assign kha = ~KHA;  //complement 
assign KHB = ~khb;  //complement 
assign kia = ~KIA;  //complement 
assign khc = ~KHC;  //complement 
assign mdk = ~MDK;  //complement 
assign CDK =  BAD & ADD  ; 
assign cdk = ~CDK;  //complement 
assign CDL =  BAD & ADF  ; 
assign cdl = ~CDL;  //complement 
assign CDM =  BAD & ADH  ; 
assign cdm = ~CDM;  //complement 
assign CXC =  BBH & ACD  ; 
assign cxc = ~CXC;  //complement 
assign CXD =  BBH & ACF  ; 
assign cxd = ~CXD;  //complement 
assign CXE =  BBH & ACH  ; 
assign cxe = ~CXE;  //complement 
assign KIB = ~kib;  //complement 
assign kja = ~KJA;  //complement 
assign KJB = ~kjb;  //complement 
assign kka = ~KKA;  //complement 
assign NFB = ~nfb;  //complement 
assign CDN =  BAD & ADJ  ; 
assign cdn = ~CDN;  //complement 
assign CDO =  BAD & ADL  ; 
assign cdo = ~CDO;  //complement 
assign CEA =  BAE & ACA  ; 
assign cea = ~CEA;  //complement 
assign CYA =  BBI & ACA  ; 
assign cya = ~CYA;  //complement 
assign CYB =  BBI & ACC  ; 
assign cyb = ~CYB;  //complement 
assign CYC =  BBI & ACE  ; 
assign cyc = ~CYC;  //complement 
assign KKB = ~kkb;  //complement 
assign kla = ~KLA;  //complement 
assign KLB = ~klb;  //complement 
assign kma = ~KMA;  //complement 
assign NFC = ~nfc;  //complement 
assign CEB =  BAE & ACC  ; 
assign ceb = ~CEB;  //complement 
assign CEC =  BAE & ACE  ; 
assign cec = ~CEC;  //complement 
assign CED =  BAE & ACG  ; 
assign ced = ~CED;  //complement 
assign CYD =  BBI & ACG  ; 
assign cyd = ~CYD;  //complement 
assign CZA =  BBJ & ACQ  ; 
assign cza = ~CZA;  //complement 
assign CZB =  BBJ & ACB  ; 
assign czb = ~CZB;  //complement 
assign KMB = ~kmb;  //complement 
assign kna = ~KNA;  //complement 
assign KNB = ~knb;  //complement 
assign koa = ~KOA;  //complement 
assign NFD = ~nfd;  //complement 
assign CEE =  BAE & ACI  ; 
assign cee = ~CEE;  //complement 
assign CEF =  BAE & ACK  ; 
assign cef = ~CEF;  //complement 
assign CEG =  BAE & ACM  ; 
assign ceg = ~CEG;  //complement 
assign CZC =  BBJ & ACD  ; 
assign czc = ~CZC;  //complement 
assign CZD =  BBJ & ACF  ; 
assign czd = ~CZD;  //complement 
assign DAA =  BBK & ACA  ; 
assign daa = ~DAA;  //complement 
assign kob = ~KOB;  //complement 
assign kpa = ~KPA;  //complement 
assign kpb = ~KPB;  //complement 
assign kqa = ~KQA;  //complement 
assign dqq = ~DQQ;  //complement 
assign CEH =  BAE & ACO  ; 
assign ceh = ~CEH;  //complement 
assign CEI =  BAE & ADA  ; 
assign cei = ~CEI;  //complement 
assign CEJ =  BAE & ADC  ; 
assign cej = ~CEJ;  //complement 
assign DAB =  BBK & ACC  ; 
assign dab = ~DAB;  //complement 
assign DAC =  BBK & ACE  ; 
assign dac = ~DAC;  //complement 
assign DBA =  BBL & ACQ  ; 
assign dba = ~DBA;  //complement 
assign kqb = ~KQB;  //complement 
assign kra = ~KRA;  //complement 
assign krb = ~KRB;  //complement 
assign ksa = ~KSA;  //complement 
assign mdj = ~MDJ;  //complement 
assign NFG = ~nfg;  //complement 
assign NFH = ~nfh;  //complement 
assign NFI = ~nfi;  //complement 
assign gka = ~GKA;  //complement 
assign GKB = ~gkb;  //complement 
assign NFJ = ~nfj;  //complement 
assign PAK = ~pak;  //complement 
assign OIB = ~oib;  //complement 
assign OKB = ~okb;  //complement 
assign OMB = ~omb;  //complement 
assign OOB = ~oob;  //complement 
assign gkc = ~GKC;  //complement 
assign GKD = ~gkd;  //complement 
assign HTB =  GTA & GUB  ; 
assign htb = ~HTB;  //complement 
assign PAM =  PAL & PAI  ; 
assign pam = ~PAM;  //complement 
assign dki = ~DKI;  //complement 
assign HOA =  GOA & gpb & goc  |  goa & GPB & goc  |  goa & gpb & GOC  |  GOA & GPB & GOC  ; 
assign hoa = ~HOA; //complement 
assign hob =  GOA & gpb & goc  |  goa & GPB & goc  |  goa & gpb & GOC  |  goa & gpb & goc  ; 
assign HOB = ~hob;  //complement 
assign gla = ~GLA;  //complement 
assign GLB = ~glb;  //complement 
assign HRA =  GRA & gsb & grc  |  gra & GSB & grc  |  gra & gsb & GRC  |  GRA & GSB & GRC  ; 
assign hra = ~HRA; //complement 
assign hrb =  GRA & gsb & grc  |  gra & GSB & grc  |  gra & gsb & GRC  |  gra & gsb & grc  ; 
assign HRB = ~hrb;  //complement 
assign HTA =  GTA & gub  |  gta & GUB  ; 
assign hta = ~HTA;  //complement 
assign HUA =  GUA & gvb  |  gua & GVB  ; 
assign hua = ~HUA;  //complement 
assign gma = ~GMA;  //complement 
assign GMB = ~gmb;  //complement 
assign HUB =  GUA & GVB  ; 
assign hub = ~HUB;  //complement 
assign HVB =  GVA & GWB  ; 
assign hvb = ~HVB;  //complement 
assign HWB =  GWA & GXB  ; 
assign hwb = ~HWB;  //complement 
assign HVA =  GVA & gwb  |  gva & GWB  ; 
assign hva = ~HVA;  //complement 
assign HWA =  GWA & gxb  |  gwa & GXB  ; 
assign hwa = ~HWA;  //complement 
assign gna = ~GNA;  //complement 
assign GNB = ~gnb;  //complement 
assign HZA =  GZA & gze  |  gza & GZE  ; 
assign hza = ~HZA;  //complement 
assign OII = ~oii;  //complement 
assign OKI = ~oki;  //complement 
assign OMI = ~omi;  //complement 
assign OOI = ~ooi;  //complement 
assign nqb =  nai  ; 
assign NQB = ~nqb;  //complement 
assign nsb =  nba  ; 
assign NSB = ~nsb;  //complement 
assign HZB =  GZA & GZE  ; 
assign hzb = ~HZB;  //complement 
assign goa = ~GOA;  //complement 
assign GOB = ~gob;  //complement 
assign NQC =  NAI & NAJ  |  NEJ  ; 
assign nqc = ~NQC;  //complement 
assign NQD =  NAI & NAJ & NAK  |  NAK & NEJ  |  NEK  ; 
assign nqd = ~NQD; //complement 
assign NFE = ~nfe;  //complement 
assign NFF = ~nff;  //complement 
assign NPD =  NAE & NAF & NAG  |  NAG & NEF  |  NEG  ; 
assign npd = ~NPD; //complement 
assign NPC =  NAE & NAF  |  NEF  ; 
assign npc = ~NPC;  //complement 
assign gpa = ~GPA;  //complement 
assign GPB = ~gpb;  //complement 
assign gqa = ~GQA;  //complement 
assign GQB = ~gqb;  //complement 
assign dmg = ~DMG;  //complement 
assign DMH = ~dmh;  //complement 
assign OIJ = ~oij;  //complement 
assign OKJ = ~okj;  //complement 
assign OMJ = ~omj;  //complement 
assign OOJ = ~ooj;  //complement 
assign EJA =  DIB & did & dif  |  dib & DID & dif  |  dib & did & DIF  |  DIB & DID & DIF  ; 
assign eja = ~EJA; //complement 
assign ejb =  DIB & did & dif  |  dib & DID & dif  |  dib & did & DIF  |  dib & did & dif  ; 
assign EJB = ~ejb;  //complement 
assign EIA =  DIA & dic & die  |  dia & DIC & die  |  dia & dic & DIE  |  DIA & DIC & DIE  ; 
assign eia = ~EIA; //complement 
assign eib =  DIA & dic & die  |  dia & DIC & die  |  dia & dic & DIE  |  dia & dic & die  ; 
assign EIB = ~eib;  //complement 
assign dmi = ~DMI;  //complement 
assign DMJ = ~dmj;  //complement 
assign OIC = ~oic;  //complement 
assign OKC = ~okc;  //complement 
assign OMC = ~omc;  //complement 
assign OOC = ~ooc;  //complement 
assign EHA =  DHB & dhd & dhf  |  dhb & DHD & dhf  |  dhb & dhd & DHF  |  DHB & DHD & DHF  ; 
assign eha = ~EHA; //complement 
assign ehb =  DHB & dhd & dhf  |  dhb & DHD & dhf  |  dhb & dhd & DHF  |  dhb & dhd & dhf  ; 
assign EHB = ~ehb;  //complement 
assign EGA =  DHA & dhc & dhe  |  dha & DHC & dhe  |  dha & dhc & DHE  |  DHA & DHC & DHE  ; 
assign ega = ~EGA; //complement 
assign egb =  DHA & dhc & dhe  |  dha & DHC & dhe  |  dha & dhc & DHE  |  dha & dhc & dhe  ; 
assign EGB = ~egb;  //complement 
assign dmk = ~DMK;  //complement 
assign DML = ~dml;  //complement 
assign HFC =  GGB & ggd  |  ggb & GGD  ; 
assign hfc = ~HFC;  //complement 
assign HAA =  GAA & gac & gae  |  gaa & GAC & gae  |  gaa & gac & GAE  |  GAA & GAC & GAE  ; 
assign haa = ~HAA; //complement 
assign hab =  GAA & gac & gae  |  gaa & GAC & gae  |  gaa & gac & GAE  |  gaa & gac & gae  ; 
assign HAB = ~hab;  //complement 
assign HBA =  GBA & gbc & gbe  |  gba & GBC & gbe  |  gba & gbc & GBE  |  GBA & GBC & GBE  ; 
assign hba = ~HBA; //complement 
assign hbb =  GBA & gbc & gbe  |  gba & GBC & gbe  |  gba & gbc & GBE  |  gba & gbc & gbe  ; 
assign HBB = ~hbb;  //complement 
assign dna = ~DNA;  //complement 
assign DNB = ~dnb;  //complement 
assign HFD = GGD & GGB ; 
assign hfd = ~HFD ; //complement 
assign HCA =  GCA & gcc & gce  |  gca & GCC & gce  |  gca & gcc & GCE  |  GCA & GCC & GCE  ; 
assign hca = ~HCA; //complement 
assign hcb =  GCA & gcc & gce  |  gca & GCC & gce  |  gca & gcc & GCE  |  gca & gcc & gce  ; 
assign HCB = ~hcb;  //complement 
assign HDA =  GDA & gdc & gde  |  gda & GDC & gde  |  gda & gdc & GDE  |  GDA & GDC & GDE  ; 
assign hda = ~HDA; //complement 
assign hdb =  GDA & gdc & gde  |  gda & GDC & gde  |  gda & gdc & GDE  |  gda & gdc & gde  ; 
assign HDB = ~hdb;  //complement 
assign dnc = ~DNC;  //complement 
assign DND = ~dnd;  //complement 
assign HHC =  GIB & gid  |  gib & GID  ; 
assign hhc = ~HHC;  //complement 
assign HEA =  GEA & gec & gfb  |  gea & GEC & gfb  |  gea & gec & GFB  |  GEA & GEC & GFB  ; 
assign hea = ~HEA; //complement 
assign heb =  GEA & gec & gfb  |  gea & GEC & gfb  |  gea & gec & GFB  |  gea & gec & gfb  ; 
assign HEB = ~heb;  //complement 
assign HFA =  GFA & gfc & gfe  |  gfa & GFC & gfe  |  gfa & gfc & GFE  |  GFA & GFC & GFE  ; 
assign hfa = ~HFA; //complement 
assign hfb =  GFA & gfc & gfe  |  gfa & GFC & gfe  |  gfa & gfc & GFE  |  gfa & gfc & gfe  ; 
assign HFB = ~hfb;  //complement 
assign dne = ~DNE;  //complement 
assign DNF = ~dnf;  //complement 
assign HHD = GID & GIB ; 
assign hhd = ~HHD ; //complement 
assign HGA =  GGA & ggc & ghb  |  gga & GGC & ghb  |  gga & ggc & GHB  |  GGA & GGC & GHB  ; 
assign hga = ~HGA; //complement 
assign hgb =  GGA & ggc & ghb  |  gga & GGC & ghb  |  gga & ggc & GHB  |  gga & ggc & ghb  ; 
assign HGB = ~hgb;  //complement 
assign HHA =  GHA & ghc & ghe  |  gha & GHC & ghe  |  gha & ghc & GHE  |  GHA & GHC & GHE  ; 
assign hha = ~HHA; //complement 
assign hhb =  GHA & ghc & ghe  |  gha & GHC & ghe  |  gha & ghc & GHE  |  gha & ghc & ghe  ; 
assign HHB = ~hhb;  //complement 
assign dng = ~DNG;  //complement 
assign DNH = ~dnh;  //complement 
assign jna = ~JNA;  //complement 
assign HIA =  GIA & gic & gjb  |  gia & GIC & gjb  |  gia & gic & GJB  |  GIA & GIC & GJB  ; 
assign hia = ~HIA; //complement 
assign hib =  GIA & gic & gjb  |  gia & GIC & gjb  |  gia & gic & GJB  |  gia & gic & gjb  ; 
assign HIB = ~hib;  //complement 
assign HJA =  GJA & gjc & gkb  |  gja & GJC & gkb  |  gja & gjc & GKB  |  GJA & GJC & GKB  ; 
assign hja = ~HJA; //complement 
assign hjb =  GJA & gjc & gkb  |  gja & GJC & gkb  |  gja & gjc & GKB  |  gja & gjc & gkb  ; 
assign HJB = ~hjb;  //complement 
assign dni = ~DNI;  //complement 
assign DNJ = ~dnj;  //complement 
assign jnb = ~JNB;  //complement 
assign HKA =  GKA & gkc & glb  |  gka & GKC & glb  |  gka & gkc & GLB  |  GKA & GKC & GLB  ; 
assign hka = ~HKA; //complement 
assign hkb =  GKA & gkc & glb  |  gka & GKC & glb  |  gka & gkc & GLB  |  gka & gkc & glb  ; 
assign HKB = ~hkb;  //complement 
assign HLA =  GLA & glc & gmb  |  gla & GLC & gmb  |  gla & glc & GMB  |  GLA & GLC & GMB  ; 
assign hla = ~HLA; //complement 
assign hlb =  GLA & glc & gmb  |  gla & GLC & gmb  |  gla & glc & GMB  |  gla & glc & gmb  ; 
assign HLB = ~hlb;  //complement 
assign CEK =  BAE & ADE  ; 
assign cek = ~CEK;  //complement 
assign CEL =  BAE & ADG  ; 
assign cel = ~CEL;  //complement 
assign CEM =  BAE & ADI  ; 
assign cem = ~CEM;  //complement 
assign DBB =  BBL & ACB  ; 
assign dbb = ~DBB;  //complement 
assign DBC =  BBL & ACD  ; 
assign dbc = ~DBC;  //complement 
assign DCA =  BBM & ACA  ; 
assign dca = ~DCA;  //complement 
assign ksb = ~KSB;  //complement 
assign kta = ~KTA;  //complement 
assign ktb = ~KTB;  //complement 
assign kua = ~KUA;  //complement 
assign gwa = ~GWA;  //complement 
assign CEN =  BAE & ADK  ; 
assign cen = ~CEN;  //complement 
assign CFA =  BAF & ACQ  ; 
assign cfa = ~CFA;  //complement 
assign CFB =  BAF & ACB  ; 
assign cfb = ~CFB;  //complement 
assign DCB =  BBM & ACC  ; 
assign dcb = ~DCB;  //complement 
assign DDA =  BBN & ACQ  ; 
assign dda = ~DDA;  //complement 
assign DDB =  BBN & ACB  ; 
assign ddb = ~DDB;  //complement 
assign kub = ~KUB;  //complement 
assign kva = ~KVA;  //complement 
assign kvb = ~KVB;  //complement 
assign kwa = ~KWA;  //complement 
assign OIK = ~oik;  //complement 
assign OKK = ~okk;  //complement 
assign OMK = ~omk;  //complement 
assign OOK = ~ook;  //complement 
assign CFC =  BAF & ACD  ; 
assign cfc = ~CFC;  //complement 
assign CFD =  BAF & ACF  ; 
assign cfd = ~CFD;  //complement 
assign CFE =  BAF & ACH  ; 
assign cfe = ~CFE;  //complement 
assign DEA =  BBO & ACA  ; 
assign dea = ~DEA;  //complement 
assign DFA =  BBP & ACQ  ; 
assign dfa = ~DFA;  //complement 
assign kwb = ~KWB;  //complement 
assign kxa = ~KXA;  //complement 
assign kxb = ~KXB;  //complement 
assign kya = ~KYA;  //complement 
assign OIE = ~oie;  //complement 
assign OKE = ~oke;  //complement 
assign OME = ~ome;  //complement 
assign OOE = ~ooe;  //complement 
assign CFF =  BAF & ACJ  ; 
assign cff = ~CFF;  //complement 
assign CFG =  BAF & ACL  ; 
assign cfg = ~CFG;  //complement 
assign CFH =  BAF & ACN  ; 
assign cfh = ~CFH;  //complement 
assign kyb = ~KYB;  //complement 
assign kza = ~KZA;  //complement 
assign kzb = ~KZB;  //complement 
assign kzc = ~KZC;  //complement 
assign NSC =  NBA & NBB  |  NFB  ; 
assign nsc = ~NSC;  //complement 
assign NSD =  NBA & NBB & NBC  |  NBC & NFB  |  NFC  ; 
assign nsd = ~NSD; //complement 
assign CFI =  BAF & ACP  ; 
assign cfi = ~CFI;  //complement 
assign CFJ =  BAF & ADB  ; 
assign cfj = ~CFJ;  //complement 
assign CFK =  BAF & ADD  ; 
assign cfk = ~CFK;  //complement 
assign kzg = ~KZG;  //complement 
assign kzi = ~KZI;  //complement 
assign pad = ~PAD;  //complement 
assign pae = ~PAE;  //complement 
assign CFL =  BAF & ADF  ; 
assign cfl = ~CFL;  //complement 
assign CFM =  BAF & ADH  ; 
assign cfm = ~CFM;  //complement 
assign CFN =  BAF & ADJ  ; 
assign cfn = ~CFN;  //complement 
assign kzj = ~KZJ;  //complement 
assign kzl = ~KZL;  //complement 
assign kzm = ~KZM;  //complement 
assign ntb = nbe; 
assign NTB = ~ntb; //complement 
assign nxb =  nae  |  naf  |  nag  |  nah  ;
assign NXB = ~nxb;  //complement 
assign CGA =  BAG & ACA  ; 
assign cga = ~CGA;  //complement 
assign CGB =  BAG & ACC  ; 
assign cgb = ~CGB;  //complement 
assign CGC =  BAG & ACE  ; 
assign cgc = ~CGC;  //complement 
assign mee = ~MEE;  //complement 
assign mef = ~MEF;  //complement 
assign pfa = ~PFA;  //complement 
assign HZC =  GZD  ; 
assign hzc = ~HZC;  //complement 
assign HEC =  GFD  ; 
assign hec = ~HEC;  //complement 
assign EFA =  DGH & dgk  |  dgh & DGK  ; 
assign efa = ~EFA;  //complement 
assign CGD =  BAG & ACG  ; 
assign cgd = ~CGD;  //complement 
assign CGE =  BAG & ACI  ; 
assign cge = ~CGE;  //complement 
assign CGF =  BAG & ACK  ; 
assign cgf = ~CGF;  //complement 
assign pfb = ~PFB;  //complement 
assign pfc = ~PFC;  //complement 
assign pfd = ~PFD;  //complement 
assign pab = ~PAB;  //complement 
assign med = ~MED;  //complement 
assign mea = ~MEA;  //complement 
assign meh = ~MEH;  //complement 
assign OID = ~oid;  //complement 
assign OKD = ~okd;  //complement 
assign OMD = ~omd;  //complement 
assign OOD = ~ood;  //complement 
assign gwb = ~GWB;  //complement 
assign npb =  nae  ; 
assign NPB = ~npb;  //complement 
assign NNB =  NFN  ; 
assign nnb = ~NNB;  //complement 
assign OIF = ~oif;  //complement 
assign OKF = ~okf;  //complement 
assign OMF = ~omf;  //complement 
assign OOF = ~oof;  //complement 
assign gra = ~GRA;  //complement 
assign GRB = ~grb;  //complement 
assign pdf = ~PDF;  //complement 
assign pdg = ~PDG;  //complement 
assign pdh = ~PDH;  //complement 
assign gsa = ~GSA;  //complement 
assign GSB = ~gsb;  //complement 
assign pdk = ~PDK;  //complement 
assign pdl = ~PDL;  //complement 
assign pdj = ~PDJ;  //complement 
assign pdn = ~PDN;  //complement 
assign gta = ~GTA;  //complement 
assign GTB = ~gtb;  //complement 
assign pdp = ~PDP;  //complement 
assign pdo = ~PDO;  //complement 
assign gua = ~GUA;  //complement 
assign GUB = ~gub;  //complement 
assign OIL = ~oil;  //complement 
assign OKL = ~okl;  //complement 
assign OML = ~oml;  //complement 
assign OOL = ~ool;  //complement 
assign HZE =  GZF & gzn  |  gzf & GZN  ; 
assign hze = ~HZE;  //complement 
assign peb = ~PEB;  //complement 
assign gva = ~GVA;  //complement 
assign GVB = ~gvb;  //complement 
assign pec = ~PEC;  //complement 
assign jzc = ~JZC;  //complement 
assign ped = ~PED;  //complement 
assign gxa = ~GXA;  //complement 
assign GXB = ~gxb;  //complement 
assign pac = ~PAC;  //complement 
assign nxc =  nai  |  naj  |  nak  |  nal  ;
assign NXC = ~nxc;  //complement 
assign nxd =  nam  |  nan  |  nao  |  nap  ;
assign NXD = ~nxd;  //complement 
assign nxe =  nba  |  nbb  |  nbc  |  nbd  ;
assign NXE = ~nxe;  //complement 
assign nxf =  nbe  |  nbf  |  nbg  |  nbh  ;
assign NXF = ~nxf;  //complement 
assign NNC =  NFM & NBN  |  NFN  ; 
assign nnc = ~NNC;  //complement 
assign jaa = ~JAA;  //complement 
assign JAB = ~jab;  //complement 
assign jba = ~JBA;  //complement 
assign JBB = ~jbb;  //complement 
assign dnk = ~DNK;  //complement 
assign DNL = ~dnl;  //complement 
assign pej = ~PEJ;  //complement 
assign HMA =  GMA & gmc & gnb  |  gma & GMC & gnb  |  gma & gmc & GNB  |  GMA & GMC & GNB  ; 
assign hma = ~HMA; //complement 
assign hmb =  GMA & gmc & gnb  |  gma & GMC & gnb  |  gma & gmc & GNB  |  gma & gmc & gnb  ; 
assign HMB = ~hmb;  //complement 
assign HNA =  GNA & gnc & gob  |  gna & GNC & gob  |  gna & gnc & GOB  |  GNA & GNC & GOB  ; 
assign hna = ~HNA; //complement 
assign hnb =  GNA & gnc & gob  |  gna & GNC & gob  |  gna & gnc & GOB  |  gna & gnc & gob  ; 
assign HNB = ~hnb;  //complement 
assign doa = ~DOA;  //complement 
assign DOB = ~dob;  //complement 
assign pek = ~PEK;  //complement 
assign HPA =  GPA & gpc & gqb  |  gpa & GPC & gqb  |  gpa & gpc & GQB  |  GPA & GPC & GQB  ; 
assign hpa = ~HPA; //complement 
assign hpb =  GPA & gpc & gqb  |  gpa & GPC & gqb  |  gpa & gpc & GQB  |  gpa & gpc & gqb  ; 
assign HPB = ~hpb;  //complement 
assign HQA =  GQA & gqc & grb  |  gqa & GQC & grb  |  gqa & gqc & GRB  |  GQA & GQC & GRB  ; 
assign hqa = ~HQA; //complement 
assign hqb =  GQA & gqc & grb  |  gqa & GQC & grb  |  gqa & gqc & GRB  |  gqa & gqc & grb  ; 
assign HQB = ~hqb;  //complement 
assign doc = ~DOC;  //complement 
assign DOD = ~dod;  //complement 
assign pep = ~PEP;  //complement 
assign HSA =  GSA & gsc & gtb  |  gsa & GSC & gtb  |  gsa & gsc & GTB  |  GSA & GSC & GTB  ; 
assign hsa = ~HSA; //complement 
assign hsb =  GSA & gsc & gtb  |  gsa & GSC & gtb  |  gsa & gsc & GTB  |  gsa & gsc & gtb  ; 
assign HSB = ~hsb;  //complement 
assign LZC =  ZZO  ; 
assign lzc = ~LZC;  //complement 
assign LED =  KEA & KFB  ; 
assign led = ~LED;  //complement 
assign LDB =  JDA & JEB  ; 
assign ldb = ~LDB;  //complement 
assign doe = ~DOE;  //complement 
assign DOF = ~dof;  //complement 
assign pel = ~PEL;  //complement 
assign LBA =  JBA & jbc & kba  |  jba & JBC & kba  |  jba & jbc & KBA  |  JBA & JBC & KBA  ; 
assign lba = ~LBA; //complement 
assign lbb =  JBA & jbc & kba  |  jba & JBC & kba  |  jba & jbc & KBA  |  jba & jbc & kba  ; 
assign LBB = ~lbb;  //complement 
assign LBC =  KBC & kcb & jcb  |  kbc & KCB & jcb  |  kbc & kcb & JCB  |  KBC & KCB & JCB  ; 
assign lbc = ~LBC; //complement 
assign lbd =  KBC & kcb & jcb  |  kbc & KCB & jcb  |  kbc & kcb & JCB  |  kbc & kcb & jcb  ; 
assign LBD = ~lbd;  //complement 
assign dog = ~DOG;  //complement 
assign DOH = ~doh;  //complement 
assign OIM = ~oim;  //complement 
assign OKM = ~okm;  //complement 
assign OMM = ~omm;  //complement 
assign OOM = ~oom;  //complement 
assign LCA =  JCA & jcc & kca  |  jca & JCC & kca  |  jca & jcc & KCA  |  JCA & JCC & KCA  ; 
assign lca = ~LCA; //complement 
assign lcb =  JCA & jcc & kca  |  jca & JCC & kca  |  jca & jcc & KCA  |  jca & jcc & kca  ; 
assign LCB = ~lcb;  //complement 
assign LCC =  KCA & kcc & jdb  |  kca & KCC & jdb  |  kca & kcc & JDB  |  KCA & KCC & JDB  ; 
assign lcc = ~LCC; //complement 
assign lcd =  KCA & kcc & jdb  |  kca & KCC & jdb  |  kca & kcc & JDB  |  kca & kcc & jdb  ; 
assign LCD = ~lcd;  //complement 
assign doi = ~DOI;  //complement 
assign DOJ = ~doj;  //complement 
assign gnc = ~GNC;  //complement 
assign LDA =  JDA & jeb  |  jda & JEB  ; 
assign lda = ~LDA;  //complement 
assign LDC =  KDA & kdc & keb  |  kda & KDC & keb  |  kda & kdc & KEB  |  KDA & KDC & KEB  ; 
assign ldc = ~LDC; //complement 
assign ldd =  KDA & kdc & keb  |  kda & KDC & keb  |  kda & kdc & KEB  |  kda & kdc & keb  ; 
assign LDD = ~ldd;  //complement 
assign dok = ~DOK;  //complement 
assign DOL = ~dol;  //complement 
assign peg = ~PEG;  //complement 
assign LEA =  JEA & jec & jfb  |  jea & JEC & jfb  |  jea & jec & JFB  |  JEA & JEC & JFB  ; 
assign lea = ~LEA; //complement 
assign leb =  JEA & jec & jfb  |  jea & JEC & jfb  |  jea & jec & JFB  |  jea & jec & jfb  ; 
assign LEB = ~leb;  //complement 
assign LEC =  KEA & kfb  |  kea & KFB  ; 
assign lec = ~LEC;  //complement 
assign dom = ~DOM;  //complement 
assign DON = ~don;  //complement 
assign peh = ~PEH;  //complement 
assign LFA =  JFA & jgb & kfa  |  jfa & JGB & kfa  |  jfa & jgb & KFA  |  JFA & JGB & KFA  ; 
assign lfa = ~LFA; //complement 
assign lfb =  JFA & jgb & kfa  |  jfa & JGB & kfa  |  jfa & jgb & KFA  |  jfa & jgb & kfa  ; 
assign LFB = ~lfb;  //complement 
assign LGA =  JGA & jgc & jhb  |  jga & JGC & jhb  |  jga & jgc & JHB  |  JGA & JGC & JHB  ; 
assign lga = ~LGA; //complement 
assign lgb =  JGA & jgc & jhb  |  jga & JGC & jhb  |  jga & jgc & JHB  |  jga & jgc & jhb  ; 
assign LGB = ~lgb;  //complement 
assign CGG =  BAG & ACM  ; 
assign cgg = ~CGG;  //complement 
assign CGH =  BAG & ACO  ; 
assign cgh = ~CGH;  //complement 
assign CGI =  BAG & ADA  ; 
assign cgi = ~CGI;  //complement 
assign gae = ~GAE;  //complement 
assign naa = ~NAA;  //complement 
assign nab = ~NAB;  //complement 
assign nac = ~NAC;  //complement 
assign gsc = ~GSC;  //complement 
assign OHF = ~ohf;  //complement 
assign CGJ =  BAG & ADC  ; 
assign cgj = ~CGJ;  //complement 
assign CGK =  BAG & ADE  ; 
assign cgk = ~CGK;  //complement 
assign CGL =  BAG & ADG  ; 
assign cgl = ~CGL;  //complement 
assign oja = ~OJA;  //complement 
assign ola = ~OLA;  //complement 
assign ona = ~ONA;  //complement 
assign opa = ~OPA;  //complement 
assign nad = ~NAD;  //complement 
assign nae = ~NAE;  //complement 
assign CGM =  BAG & ADI  ; 
assign cgm = ~CGM;  //complement 
assign CHA =  BAH & ACQ  ; 
assign cha = ~CHA;  //complement 
assign CHB =  BAH & ACB  ; 
assign chb = ~CHB;  //complement 
assign naf = ~NAF;  //complement 
assign ojb = ~OJB;  //complement 
assign olb = ~OLB;  //complement 
assign onb = ~ONB;  //complement 
assign opb = ~OPB;  //complement 
assign nag = ~NAG;  //complement 
assign CHC =  BAH & ACD  ; 
assign chc = ~CHC;  //complement 
assign CHD =  BAH & ACF  ; 
assign chd = ~CHD;  //complement 
assign CHE =  BAH & ACH  ; 
assign che = ~CHE;  //complement 
assign nah = ~NAH;  //complement 
assign nai = ~NAI;  //complement 
assign naj = ~NAJ;  //complement 
assign CHF =  BAH & ACJ  ; 
assign chf = ~CHF;  //complement 
assign CHG =  BAH & ACL  ; 
assign chg = ~CHG;  //complement 
assign CHH =  BAH & ACN  ; 
assign chh = ~CHH;  //complement 
assign nak = ~NAK;  //complement 
assign nal = ~NAL;  //complement 
assign nam = ~NAM;  //complement 
assign CHI =  BAH & ACP  ; 
assign chi = ~CHI;  //complement 
assign CHJ =  BAH & ADB  ; 
assign chj = ~CHJ;  //complement 
assign CHK =  BAH & ADD  ; 
assign chk = ~CHK;  //complement 
assign nan = ~NAN;  //complement 
assign nao = ~NAO;  //complement 
assign nap = ~NAP;  //complement 
assign CHL =  BAH & ADF  ; 
assign chl = ~CHL;  //complement 
assign CHM =  BAH & ADH  ; 
assign chm = ~CHM;  //complement 
assign CIA =  BAI & ACA  ; 
assign cia = ~CIA;  //complement 
assign nbj = ~NBJ;  //complement 
assign nbk = ~NBK;  //complement 
assign NFK = ~nfk;  //complement 
assign nbl = ~NBL;  //complement 
assign NFL = ~nfl;  //complement 
assign CIB =  BAI & ACC  ; 
assign cib = ~CIB;  //complement 
assign CIC =  BAI & ACE  ; 
assign cic = ~CIC;  //complement 
assign CID =  BAI & ACG  ; 
assign cid = ~CID;  //complement 
assign nbm = ~NBM;  //complement 
assign NFM = ~nfm;  //complement 
assign nbn = ~NBN;  //complement 
assign NFN = ~nfn;  //complement 
assign nbo = ~NBO;  //complement 
assign NFO = ~nfo;  //complement 
assign nbd = ~NBD;  //complement 
assign jja = ~JJA;  //complement 
assign JJB = ~jjb;  //complement 
assign LGC =  KGA & khb  |  kga & KHB  ; 
assign lgc = ~LGC;  //complement 
assign LHA =  JHA & jib & kha  |  jha & JIB & kha  |  jha & jib & KHA  |  JHA & JIB & KHA  ; 
assign lha = ~LHA; //complement 
assign lhb =  JHA & jib & kha  |  jha & JIB & kha  |  jha & jib & KHA  |  jha & jib & kha  ; 
assign LHB = ~lhb;  //complement 
assign jca = ~JCA;  //complement 
assign JCB = ~jcb;  //complement 
assign nbf = ~NBF;  //complement 
assign LIA =  JIA & jjb & kia  |  jia & JJB & kia  |  jia & jjb & KIA  |  JIA & JJB & KIA  ; 
assign lia = ~LIA; //complement 
assign lib =  JIA & jjb & kia  |  jia & JJB & kia  |  jia & jjb & KIA  |  jia & jjb & kia  ; 
assign LIB = ~lib;  //complement 
assign LJA =  JJA & jkb & kja  |  jja & JKB & kja  |  jja & jkb & KJA  |  JJA & JKB & KJA  ; 
assign lja = ~LJA; //complement 
assign ljb =  JJA & jkb & kja  |  jja & JKB & kja  |  jja & jkb & KJA  |  jja & jkb & kja  ; 
assign LJB = ~ljb;  //complement 
assign jda = ~JDA;  //complement 
assign JDB = ~jdb;  //complement 
assign nbh = ~NBH;  //complement 
assign LKA =  JKA & jlb & kka  |  jka & JLB & kka  |  jka & jlb & KKA  |  JKA & JLB & KKA  ; 
assign lka = ~LKA; //complement 
assign lkb =  JKA & jlb & kka  |  jka & JLB & kka  |  jka & jlb & KKA  |  jka & jlb & kka  ; 
assign LKB = ~lkb;  //complement 
assign LLA =  JLA & jmb & kla  |  jla & JMB & kla  |  jla & jmb & KLA  |  JLA & JMB & KLA  ; 
assign lla = ~LLA; //complement 
assign llb =  JLA & jmb & kla  |  jla & JMB & kla  |  jla & jmb & KLA  |  jla & jmb & kla  ; 
assign LLB = ~llb;  //complement 
assign jea = ~JEA;  //complement 
assign JEB = ~jeb;  //complement 
assign NTC =  NBE & NBF  |  NFF  ; 
assign ntc = ~NTC;  //complement 
assign LMA =  JMA & jnb & kma  |  jma & JNB & kma  |  jma & jnb & KMA  |  JMA & JNB & KMA  ; 
assign lma = ~LMA; //complement 
assign lmb =  JMA & jnb & kma  |  jma & JNB & kma  |  jma & jnb & KMA  |  jma & jnb & kma  ; 
assign LMB = ~lmb;  //complement 
assign LNA =  JNA & job & kna  |  jna & JOB & kna  |  jna & job & KNA  |  JNA & JOB & KNA  ; 
assign lna = ~LNA; //complement 
assign lnb =  JNA & job & kna  |  jna & JOB & kna  |  jna & job & KNA  |  jna & job & kna  ; 
assign LNB = ~lnb;  //complement 
assign jfa = ~JFA;  //complement 
assign JFB = ~jfb;  //complement 
assign nbi = ~NBI;  //complement 
assign LOA =  JOA & jpb & koa  |  joa & JPB & koa  |  joa & jpb & KOA  |  JOA & JPB & KOA  ; 
assign loa = ~LOA; //complement 
assign lob =  JOA & jpb & koa  |  joa & JPB & koa  |  joa & jpb & KOA  |  joa & jpb & koa  ; 
assign LOB = ~lob;  //complement 
assign LPA =  JPA & jqb & kpa  |  jpa & JQB & kpa  |  jpa & jqb & KPA  |  JPA & JQB & KPA  ; 
assign lpa = ~LPA; //complement 
assign lpb =  JPA & jqb & kpa  |  jpa & JQB & kpa  |  jpa & jqb & KPA  |  jpa & jqb & kpa  ; 
assign LPB = ~lpb;  //complement 
assign jga = ~JGA;  //complement 
assign JGB = ~jgb;  //complement 
assign jha = ~JHA;  //complement 
assign JHB = ~jhb;  //complement 
assign LQA =  JQA & jrb & kqa  |  jqa & JRB & kqa  |  jqa & jrb & KQA  |  JQA & JRB & KQA  ; 
assign lqa = ~LQA; //complement 
assign lqb =  JQA & jrb & kqa  |  jqa & JRB & kqa  |  jqa & jrb & KQA  |  jqa & jrb & kqa  ; 
assign LQB = ~lqb;  //complement 
assign LRA =  JRA & jsb & kra  |  jra & JSB & kra  |  jra & jsb & KRA  |  JRA & JSB & KRA  ; 
assign lra = ~LRA; //complement 
assign lrb =  JRA & jsb & kra  |  jra & JSB & kra  |  jra & jsb & KRA  |  jra & jsb & kra  ; 
assign LRB = ~lrb;  //complement 
assign nba = ~NBA;  //complement 
assign nbb = ~NBB;  //complement 
assign LSA =  JSA & jtb & ksa  |  jsa & JTB & ksa  |  jsa & jtb & KSA  |  JSA & JTB & KSA  ; 
assign lsa = ~LSA; //complement 
assign lsb =  JSA & jtb & ksa  |  jsa & JTB & ksa  |  jsa & jtb & KSA  |  jsa & jtb & ksa  ; 
assign LSB = ~lsb;  //complement 
assign LTA =  JTA & jub & kta  |  jta & JUB & kta  |  jta & jub & KTA  |  JTA & JUB & KTA  ; 
assign lta = ~LTA; //complement 
assign ltb =  JTA & jub & kta  |  jta & JUB & kta  |  jta & jub & KTA  |  jta & jub & kta  ; 
assign LTB = ~ltb;  //complement 
assign nbc = ~NBC;  //complement 
assign LUA =  JUA & jvb & kua  |  jua & JVB & kua  |  jua & jvb & KUA  |  JUA & JVB & KUA  ; 
assign lua = ~LUA; //complement 
assign lub =  JUA & jvb & kua  |  jua & JVB & kua  |  jua & jvb & KUA  |  jua & jvb & kua  ; 
assign LUB = ~lub;  //complement 
assign jia = ~JIA;  //complement 
assign JIB = ~jib;  //complement 
assign LVA =  JVA & jwb & kva  |  jva & JWB & kva  |  jva & jwb & KVA  |  JVA & JWB & KVA  ; 
assign lva = ~LVA; //complement 
assign lvb =  JVA & jwb & kva  |  jva & JWB & kva  |  jva & jwb & KVA  |  jva & jwb & kva  ; 
assign LVB = ~lvb;  //complement 
assign dpa = ~DPA;  //complement 
assign DPB = ~dpb;  //complement 
assign mdl = ~MDL;  //complement 
assign mbo = ~MBO;  //complement 
assign mbl = ~MBL;  //complement 
assign mbi = ~MBI;  //complement 
assign MDI = ~mdi;  //complement 
assign mbp = ~MBP;  //complement 
assign mbn = ~MBN;  //complement 
assign dpc = ~DPC;  //complement 
assign DPD = ~dpd;  //complement 
assign ojc = ~OJC;  //complement 
assign olc = ~OLC;  //complement 
assign onc = ~ONC;  //complement 
assign opc = ~OPC;  //complement 
assign NHC =  NEE & NAF  |  NEF  ; 
assign nhc = ~NHC;  //complement 
assign NHD =  NEE & NAF & NAG  |  NEF & NAG  |  NEG  ; 
assign nhd = ~NHD; //complement 
assign dpe = ~DPE;  //complement 
assign DPF = ~dpf;  //complement 
assign NHE =  NEE & NAF & NAG & NAH  |  NEF & NAG & NAH  |  NEG & NAH  |  NEH  ; 
assign nhe = ~NHE;  //complement 
assign NIC =  NEI & NAJ  |  NEJ  ; 
assign nic = ~NIC;  //complement 
assign NID =  NEI & NAJ & NAK  |  NEJ & NAK  |  NEK  ; 
assign nid = ~NID; //complement 
assign dpg = ~DPG;  //complement 
assign DPH = ~dph;  //complement 
assign NIE =  NEI & NAJ & NAK & NAL  |  NEJ & NAK & NAL  |  NEK & NAL  |  NEL  ; 
assign nie = ~NIE;  //complement 
assign NJC =  NEM & NAN  |  NEN  ; 
assign njc = ~NJC;  //complement 
assign NJD =  NEM & NAN & NAO  |  NEN & NAO  |  NEO  ; 
assign njd = ~NJD; //complement 
assign dpi = ~DPI;  //complement 
assign DPJ = ~dpj;  //complement 
assign NJE =  NEM & NAN & NAO & NAP  |  NEN & NAO & NAP  |  NEO & NAP  |  NEP  ; 
assign nje = ~NJE;  //complement 
assign NKC =  NFA & NBB  |  NFB  ; 
assign nkc = ~NKC;  //complement 
assign NKD =  NFA & NBB & NBC  |  NFB & NBC  |  NFC  ; 
assign nkd = ~NKD; //complement 
assign dpk = ~DPK;  //complement 
assign DPL = ~dpl;  //complement 
assign NKE =  NFA & NBB & NBC & NBD  |  NFB & NBC & NBD  |  NFC & NBD  |  NFD  ; 
assign nke = ~NKE;  //complement 
assign NLC =  NFE & NBF  |  NFF  ; 
assign nlc = ~NLC;  //complement 
assign NLD =  NFE & NBF & NBG  |  NFF & NBG  |  NFG  ; 
assign nld = ~NLD; //complement 
assign dpm = ~DPM;  //complement 
assign DPN = ~dpn;  //complement 
assign nbp = ~NBP;  //complement 
assign NFP = ~nfp;  //complement 
assign nbe = ~NBE;  //complement 
assign NLE =  NFE & NBF & NBG & NBH  |  NFF & NBG & NBH  |  NFG & NBH  |  NFH  ; 
assign nle = ~NLE;  //complement 
assign dpo = ~DPO;  //complement 
assign DPP = ~dpp;  //complement 
assign nbg = ~NBG;  //complement 
assign ENC =  DKH & dkj  |  dkh & DKJ  ; 
assign enc = ~ENC;  //complement 
assign ojh = ~OJH;  //complement 
assign olh = ~OLH;  //complement 
assign onh = ~ONH;  //complement 
assign oph = ~OPH;  //complement 
assign CIE =  BAI & ACI  ; 
assign cie = ~CIE;  //complement 
assign CIF =  BAI & ACK  ; 
assign cif = ~CIF;  //complement 
assign CIG =  BAI & ACM  ; 
assign cig = ~CIG;  //complement 
assign jpb = ~JPB;  //complement 
assign jqa = ~JQA;  //complement 
assign jqb = ~JQB;  //complement 
assign CIH =  BAI & ACO  ; 
assign cih = ~CIH;  //complement 
assign CII =  BAI & ADA  ; 
assign cii = ~CII;  //complement 
assign CIJ =  BAI & ADC  ; 
assign cij = ~CIJ;  //complement 
assign jra = ~JRA;  //complement 
assign jrb = ~JRB;  //complement 
assign jsa = ~JSA;  //complement 
assign CIK =  BAI & ADE  ; 
assign cik = ~CIK;  //complement 
assign CIL =  BAI & ADG  ; 
assign cil = ~CIL;  //complement 
assign CJA =  BAJ & ACQ  ; 
assign cja = ~CJA;  //complement 
assign jsb = ~JSB;  //complement 
assign jta = ~JTA;  //complement 
assign jtb = ~JTB;  //complement 
assign CJB =  BAJ & ACB  ; 
assign cjb = ~CJB;  //complement 
assign CJC =  BAJ & ACD  ; 
assign cjc = ~CJC;  //complement 
assign CJD =  BAJ & ACF  ; 
assign cjd = ~CJD;  //complement 
assign jua = ~JUA;  //complement 
assign jub = ~JUB;  //complement 
assign jva = ~JVA;  //complement 
assign CJE =  BAJ & ACH  ; 
assign cje = ~CJE;  //complement 
assign CJF =  BAJ & ACJ  ; 
assign cjf = ~CJF;  //complement 
assign CJG =  BAJ & ACL  ; 
assign cjg = ~CJG;  //complement 
assign pbd = ~PBD;  //complement 
assign jvb = ~JVB;  //complement 
assign jwa = ~JWA;  //complement 
assign CJH =  BAJ & ACN  ; 
assign cjh = ~CJH;  //complement 
assign CJI =  BAJ & ACP  ; 
assign cji = ~CJI;  //complement 
assign CJJ =  BAJ & ADB  ; 
assign cjj = ~CJJ;  //complement 
assign jwb = ~JWB;  //complement 
assign jxa = ~JXA;  //complement 
assign jxb = ~JXB;  //complement 
assign CJK =  BAJ & ADD  ; 
assign cjk = ~CJK;  //complement 
assign CJL =  BAJ & ADF  ; 
assign cjl = ~CJL;  //complement 
assign CKA =  BAK & ACA  ; 
assign cka = ~CKA;  //complement 
assign NMC =  NFI & NBJ  |  NFJ  ; 
assign nmc = ~NMC;  //complement 
assign NMD =  NFI & NBJ & NBK  |  NFJ & NBK  |  NFK  ; 
assign nmd = ~NMD; //complement 
assign joa = ~JOA;  //complement 
assign CKB =  BAK & ACC  ; 
assign ckb = ~CKB;  //complement 
assign CKC =  BAK & ACE  ; 
assign ckc = ~CKC;  //complement 
assign CKD =  BAK & ACG  ; 
assign ckd = ~CKD;  //complement 
assign job = ~JOB;  //complement 
assign jpa = ~JPA;  //complement 
assign NME =  NFI & NBJ & NBK & NBL  |  NFJ & NBK & NBL  |  NFK & NBL  |  NFL  ; 
assign nme = ~NME;  //complement 
assign oji = ~OJI;  //complement 
assign oli = ~OLI;  //complement 
assign oni = ~ONI;  //complement 
assign opi = ~OPI;  //complement 
assign pbf = ~PBF;  //complement 
assign LWA =  JWA & jxb & kwa  |  jwa & JXB & kwa  |  jwa & jxb & KWA  |  JWA & JXB & KWA  ; 
assign lwa = ~LWA; //complement 
assign lwb =  JWA & jxb & kwa  |  jwa & JXB & kwa  |  jwa & jxb & KWA  |  jwa & jxb & kwa  ; 
assign LWB = ~lwb;  //complement 
assign LXA =  JXA & jyb & kxa  |  jxa & JYB & kxa  |  jxa & jyb & KXA  |  JXA & JYB & KXA  ; 
assign lxa = ~LXA; //complement 
assign lxb =  JXA & jyb & kxa  |  jxa & JYB & kxa  |  jxa & jyb & KXA  |  jxa & jyb & kxa  ; 
assign LXB = ~lxb;  //complement 
assign jka = ~JKA;  //complement 
assign JKB = ~jkb;  //complement 
assign pbg = ~PBG;  //complement 
assign LYA =  JYA & kya  |  jya & KYA  ; 
assign lya = ~LYA;  //complement 
assign LZA =  JZA & kza & jzd  |  jza & KZA & jzd  |  jza & kza & JZD  |  JZA & KZA & JZD  ; 
assign lza = ~LZA; //complement 
assign lzb =  JZA & kza & jzd  |  jza & KZA & jzd  |  jza & kza & JZD  |  jza & kza & jzd  ; 
assign LZB = ~lzb;  //complement 
assign jla = ~JLA;  //complement 
assign JLB = ~jlb;  //complement 
assign LZF =  JZE & kze  |  jze & KZE  ; 
assign lzf = ~LZF;  //complement 
assign ojd = ~OJD;  //complement 
assign old = ~OLD;  //complement 
assign ond = ~OND;  //complement 
assign opd = ~OPD;  //complement 
assign LZD =  JZC & kzc & kzf  |  jzc & KZC & kzf  |  jzc & kzc & KZF  |  JZC & KZC & KZF  ; 
assign lzd = ~LZD; //complement 
assign lze =  JZC & kzc & kzf  |  jzc & KZC & kzf  |  jzc & kzc & KZF  |  jzc & kzc & kzf  ; 
assign LZE = ~lze;  //complement 
assign jma = ~JMA;  //complement 
assign JMB = ~jmb;  //complement 
assign LZH =  JZG & kzg  |  jzg & KZG  ; 
assign lzh = ~LZH;  //complement 
assign LZI =  JZG & KZG  ; 
assign lzi = ~LZI;  //complement 
assign LGD =  KGA & KHB  ; 
assign lgd = ~LGD;  //complement 
assign NLB =  NFE  ; 
assign nlb = ~NLB;  //complement 
assign oje = ~OJE;  //complement 
assign ole = ~OLE;  //complement 
assign one = ~ONE;  //complement 
assign ope = ~OPE;  //complement 
assign NND =  NFM & NBN & NBO  |  NFN & NBO  |  NFO  ; 
assign nnd = ~NND; //complement 
assign NNE =  NFM & NBN & NBO & NBP  |  NFN & NBO & NBP  |  NFO & NBP  |  NFP  ; 
assign nne = ~NNE;  //complement 
assign LZJ =  JZI & kzi  |  jzi & KZI  ; 
assign lzj = ~LZJ;  //complement 
assign mab = ~MAB;  //complement 
assign MCB = ~mcb;  //complement 
assign LZP = KZM; 
assign lzp = ~LZP; //complement 
assign NJB = NEM; 
assign njb = ~NJB;  //complement 
assign NHB = NEE; 
assign nhb = ~NHB;  //complement 
assign pbh = ~PBH;  //complement 
assign LZL =  JZK & kzj  |  jzk & KZJ  ; 
assign lzl = ~LZL;  //complement 
assign mac = ~MAC;  //complement 
assign MCC = ~mcc;  //complement 
assign jya = ~JYA;  //complement 
assign jyb = ~JYB;  //complement 
assign dkj = ~DKJ;  //complement 
assign jze = ~JZE;  //complement 
assign jza = ~JZA;  //complement 
assign NUD =  NBI & NBJ & NBK  |  NBK & NFJ  |  NFK  ; 
assign nud = ~NUD; //complement 
assign jzd = ~JZD;  //complement 
assign mad = ~MAD;  //complement 
assign MCD = ~mcd;  //complement 
assign mae = ~MAE;  //complement 
assign MCE = ~mce;  //complement 
assign dqa = ~DQA;  //complement 
assign DQB = ~dqb;  //complement 
assign gaf = ~GAF;  //complement 
assign pfk = ~PFK;  //complement 
assign pfl = ~PFL;  //complement 
assign pfm = ~PFM;  //complement 
assign pfn = ~PFN;  //complement 
assign dqc = ~DQC;  //complement 
assign DQD = ~dqd;  //complement 
assign pbj = ~PBJ;  //complement 
assign pfo = ~PFO;  //complement 
assign pfp = ~PFP;  //complement 
assign pga = ~PGA;  //complement 
assign pgb = ~PGB;  //complement 
assign dqe = ~DQE;  //complement 
assign DQF = ~dqf;  //complement 
assign pgc = ~PGC;  //complement 
assign pgd = ~PGD;  //complement 
assign pge = ~PGE;  //complement 
assign pgf = ~PGF;  //complement 
assign pgg = ~PGG;  //complement 
assign pgh = ~PGH;  //complement 
assign dqg = ~DQG;  //complement 
assign DQH = ~dqh;  //complement 
assign pbk = ~PBK;  //complement 
assign pgi = ~PGI;  //complement 
assign pgk = ~PGK;  //complement 
assign dqi = ~DQI;  //complement 
assign DQJ = ~dqj;  //complement 
assign pgm = ~PGM;  //complement 
assign pgo = ~PGO;  //complement 
assign pbl = ~PBL;  //complement 
assign dqk = ~DQK;  //complement 
assign DQL = ~dql;  //complement 
assign pbn = ~PBN;  //complement 
assign pbo = ~PBO;  //complement 
assign pbp = ~PBP;  //complement 
assign dqm = ~DQM;  //complement 
assign DQN = ~dqn;  //complement 
assign LZM =  JZK & KZJ  ; 
assign lzm = ~LZM;  //complement 
assign NMB =  NFI  ; 
assign nmb = ~NMB;  //complement 
assign LYB =  JYA & KYA  ; 
assign lyb = ~LYB;  //complement 
assign LZN =  JZL & kzl  |  jzl & KZL  ; 
assign lzn = ~LZN;  //complement 
assign LZO =  JZL & KZL  ; 
assign lzo = ~LZO;  //complement 
assign dqo = ~DQO;  //complement 
assign DQP = ~dqp;  //complement 
assign pfe = ~PFE;  //complement 
assign pff = ~PFF;  //complement 
assign pfg = ~PFG;  //complement 
assign pfh = ~PFH;  //complement 
assign pfi = ~PFI;  //complement 
assign pfj = ~PFJ;  //complement 
assign CKE =  BAK & ACI  ; 
assign cke = ~CKE;  //complement 
assign CKF =  BAK & ACK  ; 
assign ckf = ~CKF;  //complement 
assign CKG =  BAK & ACM  ; 
assign ckg = ~CKG;  //complement 
assign HXA =  GXA & gyb  |  gxa & GYB  ; 
assign hxa = ~HXA;  //complement 
assign HXB =  GXA & GYB  ; 
assign hxb = ~HXB;  //complement 
assign HYB =  GYA & GZB  ; 
assign hyb = ~HYB;  //complement 
assign LYC =  KZB  ; 
assign lyc = ~LYC;  //complement 
assign HYA =  GYA & gzb  |  gya & GZB  ; 
assign hya = ~HYA;  //complement 
assign CKH =  BAK & ACO  ; 
assign ckh = ~CKH;  //complement 
assign CKI =  BAK & ADA  ; 
assign cki = ~CKI;  //complement 
assign CKJ =  BAK & ADC  ; 
assign ckj = ~CKJ;  //complement 
assign FEG = DST; 
assign feg = ~FEG; //complement 
assign FBG = DRS; 
assign fbg = ~FBG;  //complement 
assign EYG = DQR; 
assign eyg = ~EYG;  //complement 
assign EVE = DON; 
assign eve = ~EVE; //complement 
assign ETE = DNO; 
assign ete = ~ETE;  //complement 
assign ESE = DNM; 
assign ese = ~ESE;  //complement 
assign ELC = DJH; 
assign elc = ~ELC;  //complement 
assign EKC = DJG; 
assign ekc = ~EKC; //complement 
assign EDA = DGE; 
assign eda = ~EDA;  //complement 
assign EBA = DGC; 
assign eba = ~EBA;  //complement 
assign EAA = DGA; 
assign eaa = ~EAA;  //complement 
assign CKK =  BAK & ADE  ; 
assign ckk = ~CKK;  //complement 
assign CLA =  BAL & ACQ  ; 
assign cla = ~CLA;  //complement 
assign CLB =  BAL & ACB  ; 
assign clb = ~CLB;  //complement 
assign HIC = GJD; 
assign hic = ~HIC; //complement 
assign HJC = GKD; 
assign hjc = ~HJC;  //complement 
assign HKC = GLD; 
assign hkc = ~HKC;  //complement 
assign HLC = GMD; 
assign hlc = ~HLC;  //complement 
assign HMC = GND; 
assign hmc = ~HMC; //complement 
assign LCE = KDB; 
assign lce = ~LCE;  //complement 
assign LFD = KFC & KGB ; 
assign lfd = ~LFD ;  //complement 
assign LHC = khc & KIB ; 
assign lhc = ~LHC ; //complement 
assign LIC = khc & KJB ; 
assign lic = ~LIC ;  //complement 
assign LJC = KKB; 
assign ljc = ~LJC;  //complement 
assign LKC = KLB; 
assign lkc = ~LKC;  //complement 
assign CLC =  BAL & ACD  ; 
assign clc = ~CLC;  //complement 
assign CLD =  BAL & ACF  ; 
assign cld = ~CLD;  //complement 
assign CLE =  BAL & ACH  ; 
assign cle = ~CLE;  //complement 
assign LLC = KMB; 
assign llc = ~LLC; //complement 
assign LMC = KNB; 
assign lmc = ~LMC;  //complement 
assign LNC = KOB; 
assign lnc = ~LNC;  //complement 
assign LOC = KPB; 
assign loc = ~LOC;  //complement 
assign LPC = KQB; 
assign lpc = ~LPC; //complement 
assign LQC = KRB; 
assign lqc = ~LQC;  //complement 
assign LRC = KSB; 
assign lrc = ~LRC;  //complement 
assign LSC = KTB; 
assign lsc = ~LSC;  //complement 
assign LTC = KUB; 
assign ltc = ~LTC; //complement 
assign LUC = KVB; 
assign luc = ~LUC;  //complement 
assign LVC = KWB; 
assign lvc = ~LVC;  //complement 
assign LWC = KXB; 
assign lwc = ~LWC;  //complement 
assign CLF =  BAL & ACJ  ; 
assign clf = ~CLF;  //complement 
assign CLG =  BAL & ACL  ; 
assign clg = ~CLG;  //complement 
assign CLH =  BAL & ACN  ; 
assign clh = ~CLH;  //complement 
assign pba = ~PBA;  //complement 
assign pbb = ~PBB;  //complement 
assign pbc = ~PBC;  //complement 
assign pbe = ~PBE;  //complement 
assign pbi = ~PBI;  //complement 
assign pbm = ~PBM;  //complement 
assign pca = ~PCA;  //complement 
assign pce = ~PCE;  //complement 
assign pci = ~PCI;  //complement 
assign pcm = ~PCM;  //complement 
assign pde = ~PDE;  //complement 
assign CLI =  BAL & ACP  ; 
assign cli = ~CLI;  //complement 
assign CLJ =  BAL & ADB  ; 
assign clj = ~CLJ;  //complement 
assign CLK =  BAL & ADD  ; 
assign clk = ~CLK;  //complement 
assign pdi = ~PDI;  //complement 
assign pdm = ~PDM;  //complement 
assign pea = ~PEA;  //complement 
assign pee = ~PEE;  //complement 
assign pei = ~PEI;  //complement 
assign pem = ~PEM;  //complement 
assign grc = ~GRC;  //complement 
assign paf = ~PAF;  //complement 
assign CMA =  BAM & ACA  ; 
assign cma = ~CMA;  //complement 
assign CMB =  BAM & ACC  ; 
assign cmb = ~CMB;  //complement 
assign CMC =  BAM & ACE  ; 
assign cmc = ~CMC;  //complement 
assign pcb = ~PCB;  //complement 
assign pcc = ~PCC;  //complement 
assign pcd = ~PCD;  //complement 
assign CMD =  BAM & ACG  ; 
assign cmd = ~CMD;  //complement 
assign CME =  BAM & ACI  ; 
assign cme = ~CME;  //complement 
assign CMF =  BAM & ACK  ; 
assign cmf = ~CMF;  //complement 
assign pcf = ~PCF;  //complement 
assign pcg = ~PCG;  //complement 
assign pch = ~PCH;  //complement 
assign peo = ~PEO;  //complement 
assign pen = ~PEN;  //complement 
assign pah = ~PAH;  //complement 
assign maf = ~MAF;  //complement 
assign MCF = ~mcf;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign TEA = QAA; 
assign tea = ~TEA; //complement 
assign TEB = QAA; 
assign teb = ~TEB;  //complement 
assign TEC = QAA; 
assign tec = ~TEC;  //complement 
assign TED = QAA; 
assign ted = ~TED;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign mag = ~MAG;  //complement 
assign MCG = ~mcg;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign oed = ~OED;  //complement 
assign oee = ~OEE;  //complement 
assign oef = ~OEF;  //complement 
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign ofc = ~OFC;  //complement 
assign ofd = ~OFD;  //complement 
assign ofe = ~OFE;  //complement 
assign off = ~OFF;  //complement 
assign mah = ~MAH;  //complement 
assign MCH = ~mch;  //complement 
assign gyb = ~GYB;  //complement 
assign OHC = ~ohc;  //complement 
assign OHD = ~ohd;  //complement 
assign OHE = ~ohe;  //complement 
assign OGA = ~oga;  //complement 
assign OGB = ~ogb;  //complement 
assign OGC = ~ogc;  //complement 
assign OGD = ~ogd;  //complement 
assign OGE = ~oge;  //complement 
assign OGF = ~ogf;  //complement 
assign OHA = ~oha;  //complement 
assign OHB = ~ohb;  //complement 
assign mai = ~MAI;  //complement 
assign MCI = ~mci;  //complement 
assign OIG = ~oig;  //complement 
assign OKG = ~okg;  //complement 
assign OMG = ~omg;  //complement 
assign OOG = ~oog;  //complement 
assign qai = ~QAI;  //complement 
assign qaj = ~QAJ;  //complement 
assign qak = ~QAK;  //complement 
assign nbq = ~NBQ;  //complement 
assign TEE = QAB; 
assign tee = ~TEE; //complement 
assign TEF = QAB; 
assign tef = ~TEF;  //complement 
assign TEG = QAB; 
assign teg = ~TEG;  //complement 
assign TEH = QAB; 
assign teh = ~TEH;  //complement 
assign maj = ~MAJ;  //complement 
assign MCJ = ~mcj;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign mak = ~MAK;  //complement 
assign MCK = ~mck;  //complement 
assign pcj = ~PCJ;  //complement 
assign pck = ~PCK;  //complement 
assign pcl = ~PCL;  //complement 
assign pcn = ~PCN;  //complement 
assign pco = ~PCO;  //complement 
assign pcp = ~PCP;  //complement 
assign mal = ~MAL;  //complement 
assign MCL = ~mcl;  //complement 
assign mam = ~MAM;  //complement 
assign MCM = ~mcm;  //complement 
assign dra = ~DRA;  //complement 
assign DRB = ~drb;  //complement 
assign bag = ~BAG;  //complement 
assign bah = ~BAH;  //complement 
assign bao = ~BAO;  //complement 
assign bap = ~BAP;  //complement 
assign bbo = ~BBO;  //complement 
assign bbp = ~BBP;  //complement 
assign drc = ~DRC;  //complement 
assign DRD = ~drd;  //complement 
assign bbg = ~BBG;  //complement 
assign bbh = ~BBH;  //complement 
assign kze = ~KZE;  //complement 
assign kzf = ~KZF;  //complement 
assign nxg =  nbi  |  nbj  |  nbk  |  nbl  ;
assign NXG = ~nxg;  //complement 
assign dre = ~DRE;  //complement 
assign DRF = ~drf;  //complement 
assign nxi =  nae  |  naf  |  nag  |  nah  |  nai  ;
assign NXI = ~nxi;  //complement 
assign nxj =  naj  |  nak  |  nal  |  nam  |  nan  ;
assign NXJ = ~nxj;  //complement 
assign nxk =  nao  |  nap  |  nba  |  nbb  |  nbc  ;
assign NXK = ~nxk;  //complement 
assign drg = ~DRG;  //complement 
assign DRH = ~drh;  //complement 
assign nxl =  nbd  |  nbe  |  nbf  |  nbg  |  nbh  ;
assign NXL = ~nxl;  //complement 
assign LHD =  KIB & KHC  ; 
assign lhd = ~LHD;  //complement 
assign NIB =  NEI  ; 
assign nib = ~NIB;  //complement 
assign HZL =  GZL  ; 
assign hzl = ~HZL;  //complement 
assign ojk = ~OJK;  //complement 
assign olk = ~OLK;  //complement 
assign onk = ~ONK;  //complement 
assign opk = ~OPK;  //complement 
assign dri = ~DRI;  //complement 
assign DRJ = ~drj;  //complement 
assign ojl = ~OJL;  //complement 
assign oll = ~OLL;  //complement 
assign onl = ~ONL;  //complement 
assign opl = ~OPL;  //complement 
assign ojf = ~OJF;  //complement 
assign olf = ~OLF;  //complement 
assign onf = ~ONF;  //complement 
assign opf = ~OPF;  //complement 
assign mbm = ~MBM;  //complement 
assign drk = ~DRK;  //complement 
assign DRL = ~drl;  //complement 
assign NUC =  NBI & NBJ  |  NFJ  ; 
assign nuc = ~NUC;  //complement 
assign ojj = ~OJJ;  //complement 
assign olj = ~OLJ;  //complement 
assign onj = ~ONJ;  //complement 
assign opj = ~OPJ;  //complement 
assign drm = ~DRM;  //complement 
assign DRN = ~drn;  //complement 
assign acq = ~ACQ;  //complement 
assign pgn = ~PGN;  //complement 
assign pgp = ~PGP;  //complement 
assign dro = ~DRO;  //complement 
assign DRP = ~drp;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign EUE =  DOM & doo  |  dom & DOO  ; 
assign eue = ~EUE;  //complement 
assign meb = ~MEB;  //complement 
assign CMG =  BAM & ACM  ; 
assign cmg = ~CMG;  //complement 
assign CMH =  BAM & ACO  ; 
assign cmh = ~CMH;  //complement 
assign CMI =  BAM & ADA  ; 
assign cmi = ~CMI;  //complement 
assign gya = ~GYA;  //complement 
assign gza = ~GZA;  //complement 
assign gzb = ~GZB;  //complement 
assign CMJ =  BAM & ADC  ; 
assign cmj = ~CMJ;  //complement 
assign CNA =  BAN & ACQ  ; 
assign cna = ~CNA;  //complement 
assign CNB =  BAN & ACB  ; 
assign cnb = ~CNB;  //complement 
assign gze = ~GZE;  //complement 
assign LZG =  JZE & KZE  ; 
assign lzg = ~LZG;  //complement 
assign LZK =  JZI & KZI  ; 
assign lzk = ~LZK;  //complement 
assign mdn = ~MDN;  //complement 
assign CNC =  BAN & ACD  ; 
assign cnc = ~CNC;  //complement 
assign CND =  BAN & ACF  ; 
assign cnd = ~CND;  //complement 
assign CNE =  BAN & ACH  ; 
assign cne = ~CNE;  //complement 
assign NVC =  NBM & NBN  |  NFN  ; 
assign nvc = ~NVC;  //complement 
assign pag = ~PAG;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign CNF =  BAN & ACJ  ; 
assign cnf = ~CNF;  //complement 
assign CNG =  BAN & ACL  ; 
assign cng = ~CNG;  //complement 
assign CNH =  BAN & ACN  ; 
assign cnh = ~CNH;  //complement 
assign NVD =  NBM & NBN & NBO  |  NBO & NFN  |  NFO  ; 
assign nvd = ~NVD; //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign PAI = ~pai;  //complement 
assign CNI =  BAN & ACP  ; 
assign cni = ~CNI;  //complement 
assign CNJ =  BAN & ADB  ; 
assign cnj = ~CNJ;  //complement 
assign COA =  BAO & ACA  ; 
assign coa = ~COA;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign NRD =  NAM & NAN & NAO  |  NAO & NEN  |  NEO  ; 
assign nrd = ~NRD; //complement 
assign NRC =  NAM & NAN  |  NEN  ; 
assign nrc = ~NRC;  //complement 
assign COB =  BAO & ACC  ; 
assign cob = ~COB;  //complement 
assign COC =  BAO & ACE  ; 
assign coc = ~COC;  //complement 
assign COD =  BAO & ACG  ; 
assign cod = ~COD;  //complement 
assign pef = ~PEF;  //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign COE =  BAO & ACI  ; 
assign coe = ~COE;  //complement 
assign COF =  BAO & ACK  ; 
assign cof = ~COF;  //complement 
assign COG =  BAO & ACM  ; 
assign cog = ~COG;  //complement 
assign FFH =  DTS & DTU  ; 
assign ffh = ~FFH;  //complement 
assign EMD =  DKG & DKI  ; 
assign emd = ~EMD;  //complement 
assign EFB =  DGH & DGK  ; 
assign efb = ~EFB;  //complement 
assign EEB =  DGG & DGJ  ; 
assign eeb = ~EEB;  //complement 
assign ECB =  DGD & DGF  ; 
assign ecb = ~ECB;  //complement 
assign LXC =  KYB  ; 
assign lxc = ~LXC;  //complement 
assign maa = ~MAA;  //complement 
assign MCA = ~mca;  //complement 
assign COH =  BAO & ACO  ; 
assign coh = ~COH;  //complement 
assign COI =  BAO & ADA  ; 
assign coi = ~COI;  //complement 
assign CPA =  BAP & ACQ  ; 
assign cpa = ~CPA;  //complement 
assign pgj = ~PGJ;  //complement 
assign pgl = ~PGL;  //complement 
assign ojm = ~OJM;  //complement 
assign olm = ~OLM;  //complement 
assign onm = ~ONM;  //complement 
assign opm = ~OPM;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iff = ~IFF; //complement 
assign ifg = ~IFG; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign iha = ~IHA; //complement 
always@(posedge IZZ )
   begin 
 AAL <= IAL & teb |  AAM & TEB ; 
 AAM <= IAM & teb |  AAN & TEB ; 
 AAN <= IAN & teb |  AAO & TEB ; 
 AAO <= IAO & teb |  AAP & TEB ; 
 AAP <= IAP & teb |  ABA & TEB ; 
 MAN <=  LOA & loc & lpb  |  loa & LOC & lpb  |  loa & loc & LPB  |  LOA & LOC & LPB  ;
 mcn <=  LOA & loc & lpb  |  loa & LOC & lpb  |  loa & loc & LPB  |  loa & loc & lpb  ;
 DRQ <=  CYB & czb & daa  |  cyb & CZB & daa  |  cyb & czb & DAA  |  CYB & CZB & DAA  ;
 drr <=  CYB & czb & daa  |  cyb & CZB & daa  |  cyb & czb & DAA  |  cyb & czb & daa  ;
 NEA <= ZZO ; 
 NEB <= ZZO ; 
 NEC <= ZZO ; 
 MDM <= LZM ; 
 OJG <= IFG ; 
 OLG <= IFG ; 
 ONG <= IFG ; 
 OPG <= IFG ; 
 MAO <=  LPA & lpc & lqb  |  lpa & LPC & lqb  |  lpa & lpc & LQB  |  LPA & LPC & LQB  ;
 mco <=  LPA & lpc & lqb  |  lpa & LPC & lqb  |  lpa & lpc & LQB  |  lpa & lpc & lqb  ;
 DSA <=  CAO & cbo & ccn  |  cao & CBO & ccn  |  cao & cbo & CCN  |  CAO & CBO & CCN  ;
 dsb <=  CAO & cbo & ccn  |  cao & CBO & ccn  |  cao & cbo & CCN  |  cao & cbo & ccn  ;
 DGA <= CAA & cba |  caa & CBA ; 
 DGC <= CBA & CAA ; 
 MAP <=  LQA & lqc & lrb  |  lqa & LQC & lrb  |  lqa & lqc & LRB  |  LQA & LQC & LRB  ;
 mcp <=  LQA & lqc & lrb  |  lqa & LQC & lrb  |  lqa & lqc & LRB  |  lqa & lqc & lrb  ;
 DSC <=  CDN & cem & cfm  |  cdn & CEM & cfm  |  cdn & cem & CFM  |  CDN & CEM & CFM  ;
 dsd <=  CDN & cem & cfm  |  cdn & CEM & cfm  |  cdn & cem & CFM  |  cdn & cem & cfm  ;
 DNM <= CSA & cta |  csa & CTA ; 
 DNO <= CTA & CSA ; 
 MBA <=  LRA & lrc & lsb  |  lra & LRC & lsb  |  lra & lrc & LSB  |  LRA & LRC & LSB  ;
 mda <=  LRA & lrc & lsb  |  lra & LRC & lsb  |  lra & lrc & LSB  |  lra & lrc & lsb  ;
 DSE <=  CGL & chl & cik  |  cgl & CHL & cik  |  cgl & chl & CIK  |  CGL & CHL & CIK  ;
 dsf <=  CGL & chl & cik  |  cgl & CHL & cik  |  cgl & chl & CIK  |  cgl & chl & cik  ;
 DQR <= CZA & CYA ; 
 GZN <= ECB & EDA ; 
 MBB <=  LSA & lsc & ltb  |  lsa & LSC & ltb  |  lsa & lsc & LTB  |  LSA & LSC & LTB  ;
 mdb <=  LSA & lsc & ltb  |  lsa & LSC & ltb  |  lsa & lsc & LTB  |  lsa & lsc & ltb  ;
 MDQ <= ZZO ; 
 DSG <=  CJK & ckj & clj  |  cjk & CKJ & clj  |  cjk & ckj & CLJ  |  CJK & CKJ & CLJ  ;
 dsh <=  CJK & ckj & clj  |  cjk & CKJ & clj  |  cjk & ckj & CLJ  |  cjk & ckj & clj  ;
 GJD <= EVD & EVB ; 
 NED <= MBM & MDM ; 
 MBC <=  LTA & ltc & lub  |  lta & LTC & lub  |  lta & ltc & LUB  |  LTA & LTC & LUB  ;
 mdc <=  LTA & ltc & lub  |  lta & LTC & lub  |  lta & ltc & LUB  |  lta & ltc & lub  ;
 DSI <=  CMI & cni & coh  |  cmi & CNI & coh  |  cmi & cni & COH  |  CMI & CNI & COH  ;
 dsj <=  CMI & cni & coh  |  cmi & CNI & coh  |  cmi & cni & COH  |  cmi & cni & coh  ;
 AAA <= IAA & tea |  AAB & TEA ; 
 AAB <= IAB & tea |  AAC & TEA ; 
 AAC <= IAC & tea |  AAD & TEA ; 
 AAD <= IAD & tea |  AAE & TEA ; 
 AAE <= IAE & tea |  AAF & TEA ; 
 AAF <= IAF & tea |  AAG & TEA ; 
 MBD <=  LUA & luc & lvb  |  lua & LUC & lvb  |  lua & luc & LVB  |  LUA & LUC & LVB  ;
 mdd <=  LUA & luc & lvb  |  lua & LUC & lvb  |  lua & luc & LVB  |  lua & luc & lvb  ;
 AAG <= IAG & tea |  AAH & TEA ; 
 AAH <= IAH & tea |  AAI & TEA ; 
 AAI <= IAI & teb |  AAJ & TEB ; 
 AAJ <= IAJ & teb |  AAK & TEB ; 
 AAK <= IAK & teb |  AAL & TEB ; 
 MBE <=  LVA & lvc & lwb  |  lva & LVC & lwb  |  lva & lvc & LWB  |  LVA & LVC & LWB  ;
 mde <=  LVA & lvc & lwb  |  lva & LVC & lwb  |  lva & lvc & LWB  |  lva & lvc & lwb  ;
 DSK <=  CPH & cqg & crg  |  cph & CQG & crg  |  cph & cqg & CRG  |  CPH & CQG & CRG  ;
 dsl <=  CPH & cqg & crg  |  cph & CQG & crg  |  cph & cqg & CRG  |  cph & cqg & crg  ;
 DSM <=  CSF & ctf & cue  |  csf & CTF & cue  |  csf & ctf & CUE  |  CSF & CTF & CUE  ;
 dsn <=  CSF & ctf & cue  |  csf & CTF & cue  |  csf & ctf & CUE  |  csf & ctf & cue  ;
 DGD <=  CAB & cbb & cca  |  cab & CBB & cca  |  cab & cbb & CCA  |  CAB & CBB & CCA  ;
 dge <=  CAB & cbb & cca  |  cab & CBB & cca  |  cab & cbb & CCA  |  cab & cbb & cca  ;
 ABG <= IBG & tec |  ABH & TEC ; 
 ABH <= IBH & tec |  ABI & TEC ; 
 DGG <=  CAC & cbc & ccb  |  cac & CBC & ccb  |  cac & cbc & CCB  |  CAC & CBC & CCB  ;
 dgh <=  CAC & cbc & ccb  |  cac & CBC & ccb  |  cac & cbc & CCB  |  cac & cbc & ccb  ;
 ABI <= IBI & ted |  ABJ & TED ; 
 ABJ <= IBJ & ted |  ABK & TED ; 
 ABK <= IBK & ted |  ABL & TED ; 
 DGJ <=  CDB & cea & cfa  |  cdb & CEA & cfa  |  cdb & cea & CFA  |  CDB & CEA & CFA  ;
 dgk <=  CDB & cea & cfa  |  cdb & CEA & cfa  |  cdb & cea & CFA  |  cdb & cea & cfa  ;
 ABL <= IBL & ted |  ABM & TED ; 
 ABM <= IBM & ted |  ABN & TED ; 
 ABN <= IBN & ted |  ABO & TED ; 
 DHA <=  CAD & cbd & ccc  |  cad & CBD & ccc  |  cad & cbd & CCC  |  CAD & CBD & CCC  ;
 dhb <=  CAD & cbd & ccc  |  cad & CBD & ccc  |  cad & cbd & CCC  |  cad & cbd & ccc  ;
 ABO <= IBO & ted |  ABP & TED ; 
 ABP <= IBP & ted |  ZZO & TED ; 
 DHC <=  CDC & ceb & cfb  |  cdc & CEB & cfb  |  cdc & ceb & CFB  |  CDC & CEB & CFB  ;
 dhd <=  CDC & ceb & cfb  |  cdc & CEB & cfb  |  cdc & ceb & CFB  |  cdc & ceb & cfb  ;
 GLD <= ETD & ETB ; 
 DIA <=  CAE & cbe & ccd  |  cae & CBE & ccd  |  cae & cbe & CCD  |  CAE & CBE & CCD  ;
 dib <=  CAE & cbe & ccd  |  cae & CBE & ccd  |  cae & cbe & CCD  |  cae & cbe & ccd  ;
 DRS <= DBA ; 
 GBE <= FEF ; 
 GCE <= FEE ; 
 GDE <= FCF ; 
 DIC <=  CDD & cec & cfc  |  cdd & CEC & cfc  |  cdd & cec & CFC  |  CDD & CEC & CFC  ;
 did <=  CDD & cec & cfc  |  cdd & CEC & cfc  |  cdd & cec & CFC  |  cdd & cec & cfc  ;
 ABA <= IBA & tec |  ABB & TEC ; 
 ABB <= IBB & tec |  ABC & TEC ; 
 ABC <= IBC & tec |  ABD & TEC ; 
 DIE <=  CGB & chb & cia  |  cgb & CHB & cia  |  cgb & chb & CIA  |  CGB & CHB & CIA  ;
 dif <=  CGB & chb & cia  |  cgb & CHB & cia  |  cgb & chb & CIA  |  cgb & chb & cia  ;
 ABD <= IBD & tec |  ABE & TEC ; 
 ABE <= IBE & tec |  ABF & TEC ; 
 ABF <= IBF & tec |  ABG & TEC ; 
 BAA <= IAA & tee |  BAA & TEE ; 
 BAB <= IAB & tee |  BAB & TEE ; 
 BAC <= IAC & tee |  BAC & TEE ; 
 OAA <= PFA & TFA |  ICA & tfa ; 
 OAB <= PFB & TFA |  ICB & tfa ; 
 OAC <= PFC & TFA |  ICC & tfa ; 
 BAD <= IAD & tee |  BAD & TEE ; 
 BAE <= IAE & tee |  BAE & TEE ; 
 BAF <= IAF & tee |  BAF & TEE ; 
 OAD <= PFD & TFA |  ICD & tfa ; 
 OAE <= PFE & TFA |  ICE & tfa ; 
 OAF <= PFF & TFA |  ICF & tfa ; 
 BAI <= IAI & tef |  BAI & TEF ; 
 BAJ <= IAJ & tef |  BAJ & TEF ; 
 BAK <= IAK & tef |  BAK & TEF ; 
 OAG <= PFG & TFA |  ICG & tfa ; 
 OAH <= PFH & TFA |  ICH & tfa ; 
 BAL <= IAL & tef |  BAL & TEF ; 
 BAM <= IAM & tef |  BAM & TEF ; 
 BAN <= IAN & tef |  BAN & TEF ; 
 OAI <= PFI & TFB |  ICI & tfb ; 
 OAJ <= PFJ & TFB |  ICJ & tfb ; 
 OAK <= PFK & TFB |  ICK & tfb ; 
 BBI <= IBI & teh |  BBI & TEH ; 
 BBJ <= IBJ & teh |  BBJ & TEH ; 
 BBK <= IBK & teh |  BBK & TEH ; 
 OAL <= PFL & TFB |  ICL & tfb ; 
 OAM <= PFM & TFB |  ICM & tfb ; 
 OAN <= PFN & TFB |  ICN & tfb ; 
 BBL <= teh & IBL ; 
 BBM <= teh & IBM ; 
 BBN <= teh & IBN ; 
 OAO <= PFO & TFB |  ICO & tfb ; 
 OAP <= PFP & TFB |  ICP & tfb ; 
 DGF <= CDA ; 
 DLK <= CPA ; 
 DOO <= CVA ; 
 PAL <= NHE ; 
 OBA <= PGA & TFC |  IDA & tfc ; 
 OBB <= PGB & TFC |  IDB & tfc ; 
 OBC <= PGC & TFC |  IDC & tfc ; 
 OBE <= PGE & TFC |  IDE & tfc ; 
 OBF <= PGF & TFC |  IDF & tfc ; 
 OBG <= PGG & TFC |  IDG & tfc ; 
 OBD <= PGD & TFC |  IDD & tfc ; 
 nee <=  mbl  |  mdl  ; 
 MBF <=  LWA & lwc & lxb  |  lwa & LWC & lxb  |  lwa & lwc & LXB  |  LWA & LWC & LXB  ;
 mdf <=  LWA & lwc & lxb  |  lwa & LWC & lxb  |  lwa & lwc & LXB  |  lwa & lwc & lxb  ;
 DSO <=  CVE & cwd & cxd  |  cve & CWD & cxd  |  cve & cwd & CXD  |  CVE & CWD & CXD  ;
 dsp <=  CVE & cwd & cxd  |  cve & CWD & cxd  |  cve & cwd & CXD  |  cve & cwd & cxd  ;
 nef <=  mbk  |  mdk  ; 
 neg <=  mbj  |  mdj  ; 
 MBG <=  LXA & lxc & lyb  |  lxa & LXC & lyb  |  lxa & lxc & LYB  |  LXA & LXC & LYB  ;
 mdg <=  LXA & lxc & lyb  |  lxa & LXC & lyb  |  lxa & lxc & LYB  |  lxa & lxc & lyb  ;
 DSQ <=  CYC & czc & dab  |  cyc & CZC & dab  |  cyc & czc & DAB  |  CYC & CZC & DAB  ;
 dsr <=  CYC & czc & dab  |  cyc & CZC & dab  |  cyc & czc & DAB  |  cyc & czc & dab  ;
 DHE <= CGA & cha |  cga & CHA ; 
 NEH <= MDI ; 
 MBH <=  LYA & lyc & lzb  |  lya & LYC & lzb  |  lya & lyc & LZB  |  LYA & LYC & LZB  ;
 mdh <=  LYA & lyc & lzb  |  lya & LYC & lzb  |  lya & lyc & LZB  |  lya & lyc & lzb  ;
 DSS <=  DBB & dca & dda  |  dbb & DCA & dda  |  dbb & dca & DDA  |  DBB & DCA & DDA  ;
 dst <=  DBB & dca & dda  |  dbb & DCA & dda  |  dbb & dca & DDA  |  dbb & dca & dda  ;
 nei <=  mbh  |  mdi  ; 
 nej <=  mbg  |  mdh  ; 
 nek <=  mbf  |  mdg  ; 
 DTA <=  CAP & cbp & cco  |  cap & CBP & cco  |  cap & cbp & CCO  |  CAP & CBP & CCO  ;
 dtb <=  CAP & cbp & cco  |  cap & CBP & cco  |  cap & cbp & CCO  |  cap & cbp & cco  ;
 DTU <= DEA & dfa |  dea & DFA ; 
 DTV <= DFA & DEA ; 
 DTC <=  CDO & cen & cfn  |  cdo & CEN & cfn  |  cdo & cen & CFN  |  CDO & CEN & CFN  ;
 dtd <=  CDO & cen & cfn  |  cdo & CEN & cfn  |  cdo & cen & CFN  |  cdo & cen & cfn  ;
 DTE <=  CGM & chm & cil  |  cgm & CHM & cil  |  cgm & chm & CIL  |  CGM & CHM & CIL  ;
 dtf <=  CGM & chm & cil  |  cgm & CHM & cil  |  cgm & chm & CIL  |  cgm & chm & cil  ;
 BBD <= IBD & teg |  BBD & TEG ; 
 BBE <= IBE & teg |  BBE & TEG ; 
 BBF <= IBF & teg |  BBF & TEG ; 
 BBA <= IBA & teg |  BBA & TEG ; 
 BBB <= IBB & teg |  BBB & TEG ; 
 BBC <= IBC & teg |  BBC & TEG ; 
 DTG <=  CJL & ckk & clk  |  cjl & CKK & clk  |  cjl & ckk & CLK  |  CJL & CKK & CLK  ;
 dth <=  CJL & ckk & clk  |  cjl & CKK & clk  |  cjl & ckk & CLK  |  cjl & ckk & clk  ;
 DTI <=  CMJ & cnj & coi  |  cmj & CNJ & coi  |  cmj & cnj & COI  |  CMJ & CNJ & COI  ;
 dtj <=  CMJ & cnj & coi  |  cmj & CNJ & coi  |  cmj & cnj & COI  |  cmj & cnj & coi  ;
 DJA <=  CAF & cbf & cce  |  caf & CBF & cce  |  caf & cbf & CCE  |  CAF & CBF & CCE  ;
 djb <=  CAF & cbf & cce  |  caf & CBF & cce  |  caf & cbf & CCE  |  caf & cbf & cce  ;
 GZM <= EDA & ecb |  eda & ECB ; 
 DJC <=  CDE & ced & cfd  |  cde & CED & cfd  |  cde & ced & CFD  |  CDE & CED & CFD  ;
 djd <=  CDE & ced & cfd  |  cde & CED & cfd  |  cde & ced & CFD  |  cde & ced & cfd  ;
 nel <=  mbe  |  mdf  ; 
 DJE <=  CGC & chc & cib  |  cgc & CHC & cib  |  cgc & chc & CIB  |  CGC & CHC & CIB  ;
 djf <=  CGC & chc & cib  |  cgc & CHC & cib  |  cgc & chc & CIB  |  cgc & chc & cib  ;
 nem <=  mbd  |  mde  ; 
 DJG <=  CJB & cka & cla  |  cjb & CKA & cla  |  cjb & cka & CLA  |  CJB & CKA & CLA  ;
 djh <=  CJB & cka & cla  |  cjb & CKA & cla  |  cjb & cka & CLA  |  cjb & cka & cla  ;
 DKA <=  CAG & cbg & ccf  |  cag & CBG & ccf  |  cag & cbg & CCF  |  CAG & CBG & CCF  ;
 dkb <=  CAG & cbg & ccf  |  cag & CBG & ccf  |  cag & cbg & CCF  |  cag & cbg & ccf  ;
 DKC <=  CDF & cee & cfe  |  cdf & CEE & cfe  |  cdf & cee & CFE  |  CDF & CEE & CFE  ;
 dkd <=  CDF & cee & cfe  |  cdf & CEE & cfe  |  cdf & cee & CFE  |  cdf & cee & cfe  ;
 DKE <=  CGD & chd & cic  |  cgd & CHD & cic  |  cgd & chd & CIC  |  CGD & CHD & CIC  ;
 dkf <=  CGD & chd & cic  |  cgd & CHD & cic  |  cgd & chd & CIC  |  cgd & chd & cic  ;
 GND <= ERD & ERB ; 
 DKG <=  CJC & ckb & clb  |  cjc & CKB & clb  |  cjc & ckb & CLB  |  CJC & CKB & CLB  ;
 dkh <=  CJC & ckb & clb  |  cjc & CKB & clb  |  cjc & ckb & CLB  |  cjc & ckb & clb  ;
 GZF <= EEA ; 
 GFE <= FAF ; 
 GHE <= EXF ; 
 GOC <= EQD ; 
 GPC <= EPD ; 
 OBH <= PGH & TFC |  IDH & tfc ; 
 GQC <= EOD ; 
 GZK <= EBA ; 
 GZL <= EAA ; 
 GZH <= ECA ; 
 OBI <= PGI & TFD |  IDI & tfd ; 
 OBJ <= PGJ & TFD |  IDJ & tfd ; 
 OBK <= PGK & TFD |  IDK & tfd ; 
 OBL <= PGL & TFD |  IDL & tfd ; 
 OBM <= PGM & TFD |  IDM & tfd ; 
 OBN <= PGN & TFD |  IDN & tfd ; 
 JAC <= HBD ; 
 JBC <= HCE ; 
 JCC <= HDD ; 
 DIG <= CJA ; 
 OBO <= PGO & TFD |  IDO & tfd ; 
 OBP <= PGP & TFD |  IDP & tfd ; 
 JEC <= HFD ; 
 JGC <= HHD ; 
 JZG <= HZG ; 
 JZI <= HZI ; 
 JZK <= HZK ; 
 JZL <= HZL ; 
 neo <=  mbb  |  mdc  ; 
 GMD <= ESD & ESB ; 
 KBA <= JAA ; 
 kbb <= jab ; 
 KBC <= JAC ; 
 KCA <= JBA ; 
 kcb <= jbb ; 
 KCC <= JBC ; 
 KDA <= JCA ; 
 kdb <= jcb ; 
 nen <=  mbc  |  mdd  ; 
 AAQ <= TEB & AAA ; 
 GFC <=  FBG & fab & fad  |  fbg & FAB & fad  |  fbg & fab & FAD  |  FBG & FAB & FAD  ;
 gfd <=  FBG & fab & fad  |  fbg & FAB & fad  |  fbg & fab & FAD  |  fbg & fab & fad  ;
 GBC <=  FFG & feb & fed  |  ffg & FEB & fed  |  ffg & feb & FED  |  FFG & FEB & FED  ;
 gbd <=  FFG & feb & fed  |  ffg & FEB & fed  |  ffg & feb & FED  |  ffg & feb & fed  ;
 DTK <=  CPI & cqh & crh  |  cpi & CQH & crh  |  cpi & cqh & CRH  |  CPI & CQH & CRH  ;
 dtl <=  CPI & cqh & crh  |  cpi & CQH & crh  |  cpi & cqh & CRH  |  cpi & cqh & crh  ;
 nep <=  mba  |  mdb  ; 
 GGA <=  FAA & fac & fae  |  faa & FAC & fae  |  faa & fac & FAE  |  FAA & FAC & FAE  ;
 ggb <=  FAA & fac & fae  |  faa & FAC & fae  |  faa & fac & FAE  |  faa & fac & fae  ;
 GCA <=  FEA & fec & feg  |  fea & FEC & feg  |  fea & fec & FEG  |  FEA & FEC & FEG  ;
 gcb <=  FEA & fec & feg  |  fea & FEC & feg  |  fea & fec & FEG  |  fea & fec & feg  ;
 DTM <=  CSG & ctg & cuf  |  csg & CTG & cuf  |  csg & ctg & CUF  |  CSG & CTG & CUF  ;
 dtn <=  CSG & ctg & cuf  |  csg & CTG & cuf  |  csg & ctg & CUF  |  csg & ctg & cuf  ;
 GZD <= EFA & eeb |  efa & EEB ; 
 GGC <=  EYB & eyd & eyf  |  eyb & EYD & eyf  |  eyb & eyd & EYF  |  EYB & EYD & EYF  ;
 ggd <=  EYB & eyd & eyf  |  eyb & EYD & eyf  |  eyb & eyd & EYF  |  eyb & eyd & eyf  ;
 GCC <=  FDF & fdb & fdd  |  fdf & FDB & fdd  |  fdf & fdb & FDD  |  FDF & FDB & FDD  ;
 gcd <=  FDF & fdb & fdd  |  fdf & FDB & fdd  |  fdf & fdb & FDD  |  fdf & fdb & fdd  ;
 DTO <=  CVF & cwe & cxe  |  cvf & CWE & cxe  |  cvf & cwe & CXE  |  CVF & CWE & CXE  ;
 dtp <=  CVF & cwe & cxe  |  cvf & CWE & cxe  |  cvf & cwe & CXE  |  cvf & cwe & cxe  ;
 DHF <= CGA & CHA ; 
 GHA <=  EYA & eyc & eye  |  eya & EYC & eye  |  eya & eyc & EYE  |  EYA & EYC & EYE  ;
 ghb <=  EYA & eyc & eye  |  eya & EYC & eye  |  eya & eyc & EYE  |  eya & eyc & eye  ;
 GDA <=  FDA & fdc & fde  |  fda & FDC & fde  |  fda & fdc & FDE  |  FDA & FDC & FDE  ;
 gdb <=  FDA & fdc & fde  |  fda & FDC & fde  |  fda & fdc & FDE  |  fda & fdc & fde  ;
 DTQ <=  CYD & czd & dac  |  cyd & CZD & dac  |  cyd & czd & DAC  |  CYD & CZD & DAC  ;
 dtr <=  CYD & czd & dac  |  cyd & CZD & dac  |  cyd & czd & DAC  |  cyd & czd & dac  ;
 GHC <=  EYG & exb & exd  |  eyg & EXB & exd  |  eyg & exb & EXD  |  EYG & EXB & EXD  ;
 ghd <=  EYG & exb & exd  |  eyg & EXB & exd  |  eyg & exb & EXD  |  eyg & exb & exd  ;
 GDC <=  FDG & fcb & fcd  |  fdg & FCB & fcd  |  fdg & fcb & FCD  |  FDG & FCB & FCD  ;
 gdd <=  FDG & fcb & fcd  |  fdg & FCB & fcd  |  fdg & fcb & FCD  |  fdg & fcb & fcd  ;
 DTS <=  DBC & dcb & ddb  |  dbc & DCB & ddb  |  dbc & dcb & DDB  |  DBC & DCB & DDB  ;
 dtt <=  DBC & dcb & ddb  |  dbc & DCB & ddb  |  dbc & dcb & DDB  |  dbc & dcb & ddb  ;
 GMC <= ESB & esd |  esb & ESD ; 
 GIA <=  EXA & exc & exe  |  exa & EXC & exe  |  exa & exc & EXE  |  EXA & EXC & EXE  ;
 gib <=  EXA & exc & exe  |  exa & EXC & exe  |  exa & exc & EXE  |  exa & exc & exe  ;
 GEA <=  FCA & fcc & fce  |  fca & FCC & fce  |  fca & fcc & FCE  |  FCA & FCC & FCE  ;
 geb <=  FCA & fcc & fce  |  fca & FCC & fce  |  fca & fcc & FCE  |  fca & fcc & fce  ;
 GAA <=  FGA & fgc & fge  |  fga & FGC & fge  |  fga & fgc & FGE  |  FGA & FGC & FGE  ;
 gab <=  FGA & fgc & fge  |  fga & FGC & fge  |  fga & fgc & FGE  |  fga & fgc & fge  ;
 GEC <=  FBB & fbd & fbf  |  fbb & FBD & fbf  |  fbb & fbd & FBF  |  FBB & FBD & FBF  ;
 ged <=  FBB & fbd & fbf  |  fbb & FBD & fbf  |  fbb & fbd & FBF  |  fbb & fbd & fbf  ;
 GFA <=  FBA & fbc & fbe  |  fba & FBC & fbe  |  fba & fbc & FBE  |  FBA & FBC & FBE  ;
 gfb <=  FBA & fbc & fbe  |  fba & FBC & fbe  |  fba & fbc & FBE  |  fba & fbc & fbe  ;
 GIC <=  EWB & ewd & ewf  |  ewb & EWD & ewf  |  ewb & ewd & EWF  |  EWB & EWD & EWF  ;
 gid <=  EWB & ewd & ewf  |  ewb & EWD & ewf  |  ewb & ewd & EWF  |  ewb & ewd & ewf  ;
 GJA <=  EWA & ewc & ewe  |  ewa & EWC & ewe  |  ewa & ewc & EWE  |  EWA & EWC & EWE  ;
 gjb <=  EWA & ewc & ewe  |  ewa & EWC & ewe  |  ewa & ewc & EWE  |  ewa & ewc & ewe  ;
 GAC <=  FGG & ffb & ffd  |  fgg & FFB & ffd  |  fgg & ffb & FFD  |  FGG & FFB & FFD  ;
 gad <=  FGG & ffb & ffd  |  fgg & FFB & ffd  |  fgg & ffb & FFD  |  fgg & ffb & ffd  ;
 GBA <=  FFA & ffc & ffe  |  ffa & FFC & ffe  |  ffa & ffc & FFE  |  FFA & FFC & FFE  ;
 gbb <=  FFA & ffc & ffe  |  ffa & FFC & ffe  |  ffa & ffc & FFE  |  ffa & ffc & ffe  ;
 DLA <=  CAH & cbh & ccg  |  cah & CBH & ccg  |  cah & cbh & CCG  |  CAH & CBH & CCG  ;
 dlb <=  CAH & cbh & ccg  |  cah & CBH & ccg  |  cah & cbh & CCG  |  cah & cbh & ccg  ;
 oia <= ifa ; 
 oka <= ifa ; 
 oma <= ifa ; 
 ooa <= ifa ; 
 DLC <=  CDG & cef & cff  |  cdg & CEF & cff  |  cdg & cef & CFF  |  CDG & CEF & CFF  ;
 dld <=  CDG & cef & cff  |  cdg & CEF & cff  |  cdg & cef & CFF  |  cdg & cef & cff  ;
 nfa <=  map  |  mda  ; 
 DLE <=  CGE & che & cid  |  cge & CHE & cid  |  cge & che & CID  |  CGE & CHE & CID  ;
 dlf <=  CGE & che & cid  |  cge & CHE & cid  |  cge & che & CID  |  cge & che & cid  ;
 DLG <=  CJD & ckc & clc  |  cjd & CKC & clc  |  cjd & ckc & CLC  |  CJD & CKC & CLC  ;
 dlh <=  CJD & ckc & clc  |  cjd & CKC & clc  |  cjd & ckc & CLC  |  cjd & ckc & clc  ;
 GLC <= ETB & etd |  etb & ETD ; 
 DLI <=  CMB & cnb & coa  |  cmb & CNB & coa  |  cmb & cnb & COA  |  CMB & CNB & COA  ;
 dlj <=  CMB & cnb & coa  |  cmb & CNB & coa  |  cmb & cnb & COA  |  cmb & cnb & coa  ;
 DMA <=  CAI & cbi & cch  |  cai & CBI & cch  |  cai & cbi & CCH  |  CAI & CBI & CCH  ;
 dmb <=  CAI & cbi & cch  |  cai & CBI & cch  |  cai & cbi & CCH  |  cai & cbi & cch  ;
 MBJ <= LZD ; 
 DMC <=  CDH & ceg & cfg  |  cdh & CEG & cfg  |  cdh & ceg & CFG  |  CDH & CEG & CFG  ;
 dmd <=  CDH & ceg & cfg  |  cdh & CEG & cfg  |  cdh & ceg & CFG  |  cdh & ceg & cfg  ;
 MEC <= LDB & LDD |  ZZO & ldd ; 
 DME <=  CGF & chf & cie  |  cgf & CHF & cie  |  cgf & chf & CIE  |  CGF & CHF & CIE  ;
 dmf <=  CGF & chf & cie  |  cgf & CHF & cie  |  cgf & chf & CIE  |  cgf & chf & cie  ;
 oih <= iga ; 
 okh <= iga ; 
 omh <= iga ; 
 ooh <= iga ; 
 KDC <= JCC ; 
 KEA <= JDA ; 
 keb <= jdb ; 
 KFC <= JEC ; 
 GJC <= EVB & evd |  evb & EVD ; 
 KFA <= JEA ; 
 kfb <= jeb ; 
 KGA <= JFA ; 
 kgb <= jfb ; 
 MBK <= LZF ; 
 KHA <= JGA ; 
 khb <= jgb ; 
 KIA <= JHA ; 
 KHC <= JGC ; 
 MDK <= LZI ; 
 kib <= jhb ; 
 KJA <= JIA ; 
 kjb <= jib ; 
 KKA <= JJA ; 
 nfb <=  mao  |  mcp  ; 
 kkb <= jjb ; 
 KLA <= JKA ; 
 klb <= jkb ; 
 KMA <= JLA ; 
 nfc <=  man  |  mco  ; 
 kmb <= jlb ; 
 KNA <= JMA ; 
 knb <= jmb ; 
 KOA <= JNA ; 
 nfd <=  mam  |  mcn  ; 
 KOB <= JNB ; 
 KPA <= JOA ; 
 KPB <= JOB ; 
 KQA <= JPA ; 
 DQQ <= cza & CYA ; 
 KQB <= JPB ; 
 KRA <= JQA ; 
 KRB <= JQB ; 
 KSA <= JRA ; 
 MDJ <= LZG ; 
 nfg <=  maj  |  mck  ; 
 nfh <=  mai  |  mcj  ; 
 nfi <=  mah  |  mci  ; 
 GKA <=  EVA & evc & eve  |  eva & EVC & eve  |  eva & evc & EVE  |  EVA & EVC & EVE  ;
 gkb <=  EVA & evc & eve  |  eva & EVC & eve  |  eva & evc & EVE  |  eva & evc & eve  ;
 nfj <=  mag  |  mch  ; 
 pak <=  ned  |  nxi  |  nxj  |  nxk  |  nxl  ; 
 oib <= ifb ; 
 okb <= ifb ; 
 omb <= ifb ; 
 oob <= ifb ; 
 GKC <=  EUB & eud & euf  |  eub & EUD & euf  |  eub & eud & EUF  |  EUB & EUD & EUF  ;
 gkd <=  EUB & eud & euf  |  eub & EUD & euf  |  eub & eud & EUF  |  eub & eud & euf  ;
 DKI <= CNA & cma |  cna & CMA ; 
 GLA <=  EUA & euc & eue  |  eua & EUC & eue  |  eua & euc & EUE  |  EUA & EUC & EUE  ;
 glb <=  EUA & euc & eue  |  eua & EUC & eue  |  eua & euc & EUE  |  eua & euc & eue  ;
 GMA <=  ETA & etc & ete  |  eta & ETC & ete  |  eta & etc & ETE  |  ETA & ETC & ETE  ;
 gmb <=  ETA & etc & ete  |  eta & ETC & ete  |  eta & etc & ETE  |  eta & etc & ete  ;
 GNA <=  ESA & esc & ese  |  esa & ESC & ese  |  esa & esc & ESE  |  ESA & ESC & ESE  ;
 gnb <=  ESA & esc & ese  |  esa & ESC & ese  |  esa & esc & ESE  |  esa & esc & ese  ;
 oii <= igb ; 
 oki <= igb ; 
 omi <= igb ; 
 ooi <= igb ; 
 GOA <=  ERA & erc & eqb  |  era & ERC & eqb  |  era & erc & EQB  |  ERA & ERC & EQB  ;
 gob <=  ERA & erc & eqb  |  era & ERC & eqb  |  era & erc & EQB  |  era & erc & eqb  ;
 nfe <=  mal  |  mcm  ; 
 nff <=  mak  |  mcl  ; 
 GPA <=  EQA & eqc & epb  |  eqa & EQC & epb  |  eqa & eqc & EPB  |  EQA & EQC & EPB  ;
 gpb <=  EQA & eqc & epb  |  eqa & EQC & epb  |  eqa & eqc & EPB  |  eqa & eqc & epb  ;
 GQA <=  EPA & epc & eob  |  epa & EPC & eob  |  epa & epc & EOB  |  EPA & EPC & EOB  ;
 gqb <=  EPA & epc & eob  |  epa & EPC & eob  |  epa & epc & EOB  |  epa & epc & eob  ;
 DMG <=  CJE & ckd & cld  |  cje & CKD & cld  |  cje & ckd & CLD  |  CJE & CKD & CLD  ;
 dmh <=  CJE & ckd & cld  |  cje & CKD & cld  |  cje & ckd & CLD  |  cje & ckd & cld  ;
 oij <= igc ; 
 okj <= igc ; 
 omj <= igc ; 
 ooj <= igc ; 
 DMI <=  CMC & cnc & cob  |  cmc & CNC & cob  |  cmc & cnc & COB  |  CMC & CNC & COB  ;
 dmj <=  CMC & cnc & cob  |  cmc & CNC & cob  |  cmc & cnc & COB  |  cmc & cnc & cob  ;
 oic <= ifc ; 
 okc <= ifc ; 
 omc <= ifc ; 
 ooc <= ifc ; 
 DMK <=  CPB & cqa & cra  |  cpb & CQA & cra  |  cpb & cqa & CRA  |  CPB & CQA & CRA  ;
 dml <=  CPB & cqa & cra  |  cpb & CQA & cra  |  cpb & cqa & CRA  |  cpb & cqa & cra  ;
 DNA <=  CAJ & cbj & cci  |  caj & CBJ & cci  |  caj & cbj & CCI  |  CAJ & CBJ & CCI  ;
 dnb <=  CAJ & cbj & cci  |  caj & CBJ & cci  |  caj & cbj & CCI  |  caj & cbj & cci  ;
 DNC <=  CDI & ceh & cfh  |  cdi & CEH & cfh  |  cdi & ceh & CFH  |  CDI & CEH & CFH  ;
 dnd <=  CDI & ceh & cfh  |  cdi & CEH & cfh  |  cdi & ceh & CFH  |  cdi & ceh & cfh  ;
 DNE <=  CGG & chg & cif  |  cgg & CHG & cif  |  cgg & chg & CIF  |  CGG & CHG & CIF  ;
 dnf <=  CGG & chg & cif  |  cgg & CHG & cif  |  cgg & chg & CIF  |  cgg & chg & cif  ;
 DNG <=  CJF & cke & cle  |  cjf & CKE & cle  |  cjf & cke & CLE  |  CJF & CKE & CLE  ;
 dnh <=  CJF & cke & cle  |  cjf & CKE & cle  |  cjf & cke & CLE  |  cjf & cke & cle  ;
 JNA <= HNA & hob |  hna & HOB ; 
 DNI <=  CMD & cnd & coc  |  cmd & CND & coc  |  cmd & cnd & COC  |  CMD & CND & COC  ;
 dnj <=  CMD & cnd & coc  |  cmd & CND & coc  |  cmd & cnd & COC  |  cmd & cnd & coc  ;
 JNB <= HOB & HNA ; 
 KSB <= JRB ; 
 KTA <= JSA ; 
 KTB <= JSB ; 
 KUA <= JTA ; 
 GWA <= EJA & eib |  eja & EIB ; 
 KUB <= JTB ; 
 KVA <= JUA ; 
 KVB <= JUB ; 
 KWA <= JVA ; 
 oik <= igd ; 
 okk <= igd ; 
 omk <= igd ; 
 ook <= igd ; 
 KWB <= JVB ; 
 KXA <= JWA ; 
 KXB <= JWB ; 
 KYA <= JXA ; 
 oie <= ife ; 
 oke <= ife ; 
 ome <= ife ; 
 ooe <= ife ; 
 KYB <= JXB ; 
 KZA <= JYA ; 
 KZB <= JYB ; 
 KZC <= JZA ; 
 KZG <= JZE ; 
 KZI <= JZG ; 
 PAD <=  NED & NXB & NXC  |  NHE & NXC  |  NIE  ; 
 PAE <=  NED & NXB & NXC & NXD  |  NHE & NXC & NXD  |  NIE & NXD  |  NJE  ; 
 KZJ <= JZI ; 
 KZL <= JZK ; 
 KZM <= JZL ; 
 MEE <= LGD ; 
 MEF <= LFD ; 
 PFA <= PBA ; 
 PFB <= PBB ; 
 PFC <= PBC ; 
 PFD <= PBD ; 
 PAB <= NED ; 
 MED <= LED ; 
 MEA <= LCD ; 
 MEH <= LHD ; 
 oid <= ifd ; 
 okd <= ifd ; 
 omd <= ifd ; 
 ood <= ifd ; 
 GWB <= EIB & EJA ; 
 oif <= iff ; 
 okf <= iff ; 
 omf <= iff ; 
 oof <= iff ; 
 GRA <=  EOA & eoc & enb  |  eoa & EOC & enb  |  eoa & eoc & ENB  |  EOA & EOC & ENB  ;
 grb <=  EOA & eoc & enb  |  eoa & EOC & enb  |  eoa & eoc & ENB  |  eoa & eoc & enb  ;
 PDF <= NAF & npb |  naf & NPB ; 
 PDG <= NAG & npc |  nag & NPC ; 
 PDH <= NAH & npd |  nah & NPD ; 
 GSA <=  ENA & enc & emb  |  ena & ENC & emb  |  ena & enc & EMB  |  ENA & ENC & EMB  ;
 gsb <=  ENA & enc & emb  |  ena & ENC & emb  |  ena & enc & EMB  |  ena & enc & emb  ;
 PDK <= NAK & nqc |  nak & NQC ; 
 PDL <= NAL & nqd |  nal & NQD ; 
 PDJ <= NAJ & nqb |  naj & NQB ; 
 PDN <= NAN & nrb |  nan & NRB ; 
 GTA <=  EMA & emc & elb  |  ema & EMC & elb  |  ema & emc & ELB  |  EMA & EMC & ELB  ;
 gtb <=  EMA & emc & elb  |  ema & EMC & elb  |  ema & emc & ELB  |  ema & emc & elb  ;
 PDP <= NAP & nrd |  nap & NRD ; 
 PDO <= NAO & nrc |  nao & NRC ; 
 GUA <=  ELA & elc & ekb  |  ela & ELC & ekb  |  ela & elc & EKB  |  ELA & ELC & EKB  ;
 gub <=  ELA & elc & ekb  |  ela & ELC & ekb  |  ela & elc & EKB  |  ela & elc & ekb  ;
 oil <= ige ; 
 okl <= ige ; 
 oml <= ige ; 
 ool <= ige ; 
 PEB <= NBB & nsb |  nbb & NSB ; 
 GVA <=  EKA & ekc & ejb  |  eka & EKC & ejb  |  eka & ekc & EJB  |  EKA & EKC & EJB  ;
 gvb <=  EKA & ekc & ejb  |  eka & EKC & ejb  |  eka & ekc & EJB  |  eka & ekc & ejb  ;
 PEC <= NBC & nsc |  nbc & NSC ; 
 JZC <= HZC & hzf |  hzc & HZF ; 
 PED <= NBD & nsd |  nbd & NSD ; 
 GXA <=  EIA & eic & ehb  |  eia & EIC & ehb  |  eia & eic & EHB  |  EIA & EIC & EHB  ;
 gxb <=  EIA & eic & ehb  |  eia & EIC & ehb  |  eia & eic & EHB  |  eia & eic & ehb  ;
 PAC <=  NED & NXB  |  NHE  ; 
 JAA <=  HAA & hac & hbb  |  haa & HAC & hbb  |  haa & hac & HBB  |  HAA & HAC & HBB  ;
 jab <=  HAA & hac & hbb  |  haa & HAC & hbb  |  haa & hac & HBB  |  haa & hac & hbb  ;
 JBA <=  HBA & hbc & hcb  |  hba & HBC & hcb  |  hba & hbc & HCB  |  HBA & HBC & HCB  ;
 jbb <=  HBA & hbc & hcb  |  hba & HBC & hcb  |  hba & hbc & HCB  |  hba & hbc & hcb  ;
 DNK <=  CPC & cqb & crb  |  cpc & CQB & crb  |  cpc & cqb & CRB  |  CPC & CQB & CRB  ;
 dnl <=  CPC & cqb & crb  |  cpc & CQB & crb  |  cpc & cqb & CRB  |  cpc & cqb & crb  ;
 PEJ <= NBJ & nub |  nbj & NUB ; 
 DOA <=  CAK & cbk & ccj  |  cak & CBK & ccj  |  cak & cbk & CCJ  |  CAK & CBK & CCJ  ;
 dob <=  CAK & cbk & ccj  |  cak & CBK & ccj  |  cak & cbk & CCJ  |  cak & cbk & ccj  ;
 PEK <= NBK & nuc |  nbk & NUC ; 
 DOC <=  CDJ & cei & cfi  |  cdj & CEI & cfi  |  cdj & cei & CFI  |  CDJ & CEI & CFI  ;
 dod <=  CDJ & cei & cfi  |  cdj & CEI & cfi  |  cdj & cei & CFI  |  cdj & cei & cfi  ;
 PEP <= NBP & nvd |  nbp & NVD ; 
 DOE <=  CGH & chh & cig  |  cgh & CHH & cig  |  cgh & chh & CIG  |  CGH & CHH & CIG  ;
 dof <=  CGH & chh & cig  |  cgh & CHH & cig  |  cgh & chh & CIG  |  cgh & chh & cig  ;
 PEL <= NBL & nud |  nbl & NUD ; 
 DOG <=  CJG & ckf & clf  |  cjg & CKF & clf  |  cjg & ckf & CLF  |  CJG & CKF & CLF  ;
 doh <=  CJG & ckf & clf  |  cjg & CKF & clf  |  cjg & ckf & CLF  |  cjg & ckf & clf  ;
 oim <= igf ; 
 okm <= igf ; 
 omm <= igf ; 
 oom <= igf ; 
 DOI <=  CME & cne & cod  |  cme & CNE & cod  |  cme & cne & COD  |  CME & CNE & COD  ;
 doj <=  CME & cne & cod  |  cme & CNE & cod  |  cme & cne & COD  |  cme & cne & cod  ;
 GNC <= ERB & erd |  erb & ERD ; 
 DOK <=  CPD & cqc & crc  |  cpd & CQC & crc  |  cpd & cqc & CRC  |  CPD & CQC & CRC  ;
 dol <=  CPD & cqc & crc  |  cpd & CQC & crc  |  cpd & cqc & CRC  |  cpd & cqc & crc  ;
 PEG <= NBG & ntc |  nbg & NTC ; 
 DOM <=  CSB & ctb & cua  |  csb & CTB & cua  |  csb & ctb & CUA  |  CSB & CTB & CUA  ;
 don <=  CSB & ctb & cua  |  csb & CTB & cua  |  csb & ctb & CUA  |  csb & ctb & cua  ;
 PEH <= NBH & ntd |  nbh & NTD ; 
 GAE <= FFF & ffh |  fff & FFH ; 
 NAA <= MBP ; 
 NAB <= MBO ; 
 NAC <= MBN ; 
 GSC <= EMD ; 
 ohf <= ief ; 
 OJA <= IFA ; 
 OLA <= IFA ; 
 ONA <= IFA ; 
 OPA <= IFA ; 
 NAD <= MBM & mdm |  mbm & MDM ; 
 NAE <= MBL & mdl |  mbl & MDL ; 
 NAF <= MBK & mdk |  mbk & MDK ; 
 OJB <= IFB ; 
 OLB <= IFB ; 
 ONB <= IFB ; 
 OPB <= IFB ; 
 NAG <= MBJ & mdj |  mbj & MDJ ; 
 NAH <= MBI ; 
 NAI <= MBH ; 
 NAJ <= MBG & mdh |  mbg & MDH ; 
 NAK <= MBF & mdg |  mbf & MDG ; 
 NAL <= MBE & mdf |  mbe & MDF ; 
 NAM <= MBD & mde |  mbd & MDE ; 
 NAN <= MBC & mdd |  mbc & MDD ; 
 NAO <= MBB & mdc |  mbb & MDC ; 
 NAP <= MBA & mdb |  mba & MDB ; 
 NBJ <= MAG & mch |  mag & MCH ; 
 NBK <=  MAF & mcg & meh  |  maf & MCG & meh  |  maf & mcg & MEH  |  MAF & MCG & MEH  ;
 nfk <=  MAF & mcg & meh  |  maf & MCG & meh  |  maf & mcg & MEH  |  maf & mcg & meh  ;
 NBL <=  MAE & mcf & mee  |  mae & MCF & mee  |  mae & mcf & MEE  |  MAE & MCF & MEE  ;
 nfl <=  MAE & mcf & mee  |  mae & MCF & mee  |  mae & mcf & MEE  |  mae & mcf & mee  ;
 NBM <=  MAD & mce & mef  |  mad & MCE & mef  |  mad & mce & MEF  |  MAD & MCE & MEF  ;
 nfm <=  MAD & mce & mef  |  mad & MCE & mef  |  mad & mce & MEF  |  mad & mce & mef  ;
 NBN <=  MAC & mcd & med  |  mac & MCD & med  |  mac & mcd & MED  |  MAC & MCD & MED  ;
 nfn <=  MAC & mcd & med  |  mac & MCD & med  |  mac & mcd & MED  |  mac & mcd & med  ;
 NBO <=  MAB & mcc & meb  |  mab & MCC & meb  |  mab & mcc & MEB  |  MAB & MCC & MEB  ;
 nfo <=  MAB & mcc & meb  |  mab & MCC & meb  |  mab & mcc & MEB  |  mab & mcc & meb  ;
 NBD <= MAM & mcn |  mam & MCN ; 
 JJA <=  HJA & hjc & hkb  |  hja & HJC & hkb  |  hja & hjc & HKB  |  HJA & HJC & HKB  ;
 jjb <=  HJA & hjc & hkb  |  hja & HJC & hkb  |  hja & hjc & HKB  |  hja & hjc & hkb  ;
 JCA <=  HCA & hcd & hdb  |  hca & HCD & hdb  |  hca & hcd & HDB  |  HCA & HCD & HDB  ;
 jcb <=  HCA & hcd & hdb  |  hca & HCD & hdb  |  hca & hcd & HDB  |  hca & hcd & hdb  ;
 NBF <= MAK & mcl |  mak & MCL ; 
 JDA <=  HDA & hdc & heb  |  hda & HDC & heb  |  hda & hdc & HEB  |  HDA & HDC & HEB  ;
 jdb <=  HDA & hdc & heb  |  hda & HDC & heb  |  hda & hdc & HEB  |  hda & hdc & heb  ;
 NBH <= MAI & mcj |  mai & MCJ ; 
 JEA <=  HEA & hec & hfb  |  hea & HEC & hfb  |  hea & hec & HFB  |  HEA & HEC & HFB  ;
 jeb <=  HEA & hec & hfb  |  hea & HEC & hfb  |  hea & hec & HFB  |  hea & hec & hfb  ;
 JFA <=  HFA & hfc & hgb  |  hfa & HFC & hgb  |  hfa & hfc & HGB  |  HFA & HFC & HGB  ;
 jfb <=  HFA & hfc & hgb  |  hfa & HFC & hgb  |  hfa & hfc & HGB  |  hfa & hfc & hgb  ;
 NBI <= MAH & mci |  mah & MCI ; 
 JGA <=  HGA & hgc & hhb  |  hga & HGC & hhb  |  hga & hgc & HHB  |  HGA & HGC & HHB  ;
 jgb <=  HGA & hgc & hhb  |  hga & HGC & hhb  |  hga & hgc & HHB  |  hga & hgc & hhb  ;
 JHA <=  HHA & hhc & hib  |  hha & HHC & hib  |  hha & hhc & HIB  |  HHA & HHC & HIB  ;
 jhb <=  HHA & hhc & hib  |  hha & HHC & hib  |  hha & hhc & HIB  |  hha & hhc & hib  ;
 NBA <= MAP & mda |  map & MDA ; 
 NBB <= MAO & mcp |  mao & MCP ; 
 NBC <= MAN & mco |  man & MCO ; 
 JIA <=  HIA & hic & hjb  |  hia & HIC & hjb  |  hia & hic & HJB  |  HIA & HIC & HJB  ;
 jib <=  HIA & hic & hjb  |  hia & HIC & hjb  |  hia & hic & HJB  |  hia & hic & hjb  ;
 DPA <=  CAL & cbl & cck  |  cal & CBL & cck  |  cal & cbl & CCK  |  CAL & CBL & CCK  ;
 dpb <=  CAL & cbl & cck  |  cal & CBL & cck  |  cal & cbl & CCK  |  cal & cbl & cck  ;
 MDL <= LZK ; 
 MBO <= LZN ; 
 MBL <= LZH ; 
 MBI <=  LZA & lzc & lze  |  lza & LZC & lze  |  lza & lzc & LZE  |  LZA & LZC & LZE  ;
 mdi <=  LZA & lzc & lze  |  lza & LZC & lze  |  lza & lzc & LZE  |  lza & lzc & lze  ;
 MBP <= LZP ; 
 MBN <= LZL ; 
 DPC <=  CDK & cej & cfj  |  cdk & CEJ & cfj  |  cdk & cej & CFJ  |  CDK & CEJ & CFJ  ;
 dpd <=  CDK & cej & cfj  |  cdk & CEJ & cfj  |  cdk & cej & CFJ  |  cdk & cej & cfj  ;
 OJC <= IFC ; 
 OLC <= IFC ; 
 ONC <= IFC ; 
 OPC <= IFC ; 
 DPE <=  CGI & chi & cih  |  cgi & CHI & cih  |  cgi & chi & CIH  |  CGI & CHI & CIH  ;
 dpf <=  CGI & chi & cih  |  cgi & CHI & cih  |  cgi & chi & CIH  |  cgi & chi & cih  ;
 DPG <=  CJH & ckg & clg  |  cjh & CKG & clg  |  cjh & ckg & CLG  |  CJH & CKG & CLG  ;
 dph <=  CJH & ckg & clg  |  cjh & CKG & clg  |  cjh & ckg & CLG  |  cjh & ckg & clg  ;
 DPI <=  CMF & cnf & coe  |  cmf & CNF & coe  |  cmf & cnf & COE  |  CMF & CNF & COE  ;
 dpj <=  CMF & cnf & coe  |  cmf & CNF & coe  |  cmf & cnf & COE  |  cmf & cnf & coe  ;
 DPK <=  CPE & cqd & crd  |  cpe & CQD & crd  |  cpe & cqd & CRD  |  CPE & CQD & CRD  ;
 dpl <=  CPE & cqd & crd  |  cpe & CQD & crd  |  cpe & cqd & CRD  |  cpe & cqd & crd  ;
 DPM <=  CSC & ctc & cub  |  csc & CTC & cub  |  csc & ctc & CUB  |  CSC & CTC & CUB  ;
 dpn <=  CSC & ctc & cub  |  csc & CTC & cub  |  csc & ctc & CUB  |  csc & ctc & cub  ;
 NBP <=  MAA & mcb & mea  |  maa & MCB & mea  |  maa & mcb & MEA  |  MAA & MCB & MEA  ;
 nfp <=  MAA & mcb & mea  |  maa & MCB & mea  |  maa & mcb & MEA  |  maa & mcb & mea  ;
 NBE <= MAL & mcm |  mal & MCM ; 
 DPO <=  CVB & cwa & cxa  |  cvb & CWA & cxa  |  cvb & cwa & CXA  |  CVB & CWA & CXA  ;
 dpp <=  CVB & cwa & cxa  |  cvb & CWA & cxa  |  cvb & cwa & CXA  |  cvb & cwa & cxa  ;
 NBG <= MAJ & mck |  maj & MCK ; 
 OJH <= IGA ; 
 OLH <= IGA ; 
 ONH <= IGA ; 
 OPH <= IGA ; 
 JPB <= HQB & HPA ; 
 JQA <= HQA & hrb |  hqa & HRB ; 
 JQB <= HRB & HQA ; 
 JRA <= HRA & hsb |  hra & HSB ; 
 JRB <= HSB & HRA ; 
 JSA <= HSA & htb |  hsa & HTB ; 
 JSB <= HTB & HSA ; 
 JTA <= HTA & hub |  hta & HUB ; 
 JTB <= HUB & HTA ; 
 JUA <= HUA & hvb |  hua & HVB ; 
 JUB <= HVB & HUA ; 
 JVA <= HVA & hwb |  hva & HWB ; 
 PBD <= NAD ; 
 JVB <= HWB & HVA ; 
 JWA <= HWA & hxb |  hwa & HXB ; 
 JWB <= HXB & HWA ; 
 JXA <= HXA & hyb |  hxa & HYB ; 
 JXB <= HYB & HXA ; 
 JOA <= HOA & hpb |  hoa & HPB ; 
 JOB <= HPB & HOA ; 
 JPA <= HPA & hqb |  hpa & HQB ; 
 OJI <= IGB ; 
 OLI <= IGB ; 
 ONI <= IGB ; 
 OPI <= IGB ; 
 PBF <= NAF & nhb |  naf & NHB ; 
 JKA <=  HKA & hkc & hlb  |  hka & HKC & hlb  |  hka & hkc & HLB  |  HKA & HKC & HLB  ;
 jkb <=  HKA & hkc & hlb  |  hka & HKC & hlb  |  hka & hkc & HLB  |  hka & hkc & hlb  ;
 PBG <= NAG & nhc |  nag & NHC ; 
 JLA <=  HLA & hlc & hmb  |  hla & HLC & hmb  |  hla & hlc & HMB  |  HLA & HLC & HMB  ;
 jlb <=  HLA & hlc & hmb  |  hla & HLC & hmb  |  hla & hlc & HMB  |  hla & hlc & hmb  ;
 OJD <= IFD ; 
 OLD <= IFD ; 
 OND <= IFD ; 
 OPD <= IFD ; 
 JMA <=  HMA & hmc & hnb  |  hma & HMC & hnb  |  hma & hmc & HNB  |  HMA & HMC & HNB  ;
 jmb <=  HMA & hmc & hnb  |  hma & HMC & hnb  |  hma & hmc & HNB  |  hma & hmc & hnb  ;
 OJE <= IFE ; 
 OLE <= IFE ; 
 ONE <= IFE ; 
 OPE <= IFE ; 
 MAB <=  LCA & lcc & lce  |  lca & LCC & lce  |  lca & lcc & LCE  |  LCA & LCC & LCE  ;
 mcb <=  LCA & lcc & lce  |  lca & LCC & lce  |  lca & lcc & LCE  |  lca & lcc & lce  ;
 PBH <= NAH & nhd |  nah & NHD ; 
 MAC <=  LDA & ldc & leb  |  lda & LDC & leb  |  lda & ldc & LEB  |  LDA & LDC & LEB  ;
 mcc <=  LDA & ldc & leb  |  lda & LDC & leb  |  lda & ldc & LEB  |  lda & ldc & leb  ;
 JYA <= HYA & hzb |  hya & HZB ; 
 JYB <= HZB & HYA ; 
 DKJ <= CMA & CNA ; 
 JZE <= HZE ; 
 JZA <= HZA ; 
 JZD <= HZF & HZC ; 
 MAD <=  LEA & lec & lfb  |  lea & LEC & lfb  |  lea & lec & LFB  |  LEA & LEC & LFB  ;
 mcd <=  LEA & lec & lfb  |  lea & LEC & lfb  |  lea & lec & LFB  |  lea & lec & lfb  ;
 MAE <=  LFA & lfc & lgb  |  lfa & LFC & lgb  |  lfa & lfc & LGB  |  LFA & LFC & LGB  ;
 mce <=  LFA & lfc & lgb  |  lfa & LFC & lgb  |  lfa & lfc & LGB  |  lfa & lfc & lgb  ;
 DQA <=  CAM & cbm & ccl  |  cam & CBM & ccl  |  cam & cbm & CCL  |  CAM & CBM & CCL  ;
 dqb <=  CAM & cbm & ccl  |  cam & CBM & ccl  |  cam & cbm & CCL  |  cam & cbm & ccl  ;
 GAF <= FFH & FFF ; 
 PFK <= PDK & PAC |  PBK & pac ; 
 PFL <= PDL & PAC |  PBL & pac ; 
 PFM <= PDM & PAD |  PBM & pad ; 
 PFN <= PDN & PAD |  PBN & pad ; 
 DQC <=  CDL & cek & cfk  |  cdl & CEK & cfk  |  cdl & cek & CFK  |  CDL & CEK & CFK  ;
 dqd <=  CDL & cek & cfk  |  cdl & CEK & cfk  |  cdl & cek & CFK  |  cdl & cek & cfk  ;
 PBJ <= NAJ & nib |  naj & NIB ; 
 PFO <= PDO & PAD |  PBO & pad ; 
 PFP <= PDP & PAD |  PBP & pad ; 
 PGA <= PEA & PAE |  PCA & pae ; 
 PGB <= PEB & PAE |  PCB & pae ; 
 DQE <=  CGJ & chj & cii  |  cgj & CHJ & cii  |  cgj & chj & CII  |  CGJ & CHJ & CII  ;
 dqf <=  CGJ & chj & cii  |  cgj & CHJ & cii  |  cgj & chj & CII  |  cgj & chj & cii  ;
 PGC <= PEC & PAE |  PCC & pae ; 
 PGD <= PED & PAE |  PCD & pae ; 
 PGE <= PEE & PAF |  PCE & paf ; 
 PGF <= PEF & PAF |  PCF & paf ; 
 PGG <= PEG & PAF |  PCG & paf ; 
 PGH <= PEH & PAF |  PCH & paf ; 
 DQG <=  CJI & ckh & clh  |  cji & CKH & clh  |  cji & ckh & CLH  |  CJI & CKH & CLH  ;
 dqh <=  CJI & ckh & clh  |  cji & CKH & clh  |  cji & ckh & CLH  |  cji & ckh & clh  ;
 PBK <= NAK & nic |  nak & NIC ; 
 PGI <=  PCI & pag & pak  |  PEI & PAG  |  PEI & PAK  ; 
 PGK <=  PCK & pag & pak  |  PEK & PAG  |  PEK & PAK  ; 
 DQI <=  CMG & cng & cof  |  cmg & CNG & cof  |  cmg & cng & COF  |  CMG & CNG & COF  ;
 dqj <=  CMG & cng & cof  |  cmg & CNG & cof  |  cmg & cng & COF  |  cmg & cng & cof  ;
 PGM <=  PCM & pah & pam  |  PEM & PAH  |  PEM & PAM  ; 
 PGO <=  PCO & pah & pam  |  PEO & PAH  |  PEO & PAM  ; 
 PBL <= NAL & nid |  nal & NID ; 
 DQK <=  CPF & cqe & cre  |  cpf & CQE & cre  |  cpf & cqe & CRE  |  CPF & CQE & CRE  ;
 dql <=  CPF & cqe & cre  |  cpf & CQE & cre  |  cpf & cqe & CRE  |  cpf & cqe & cre  ;
 PBN <= NAN & njb |  nan & NJB ; 
 PBO <= NAO & njc |  nao & NJC ; 
 PBP <= NAP & njd |  nap & NJD ; 
 DQM <=  CSD & ctd & cuc  |  csd & CTD & cuc  |  csd & ctd & CUC  |  CSD & CTD & CUC  ;
 dqn <=  CSD & ctd & cuc  |  csd & CTD & cuc  |  csd & ctd & CUC  |  csd & ctd & cuc  ;
 DQO <=  CVC & cwb & cxb  |  cvc & CWB & cxb  |  cvc & cwb & CXB  |  CVC & CWB & CXB  ;
 dqp <=  CVC & cwb & cxb  |  cvc & CWB & cxb  |  cvc & cwb & CXB  |  cvc & cwb & cxb  ;
 PFE <= PDE & PAB |  PBE & pab ; 
 PFF <= PDF & PAB |  PBF & pab ; 
 PFG <= PDG & PAB |  PBG & pab ; 
 PFH <= PDH & PAB |  PBH & pab ; 
 PFI <= PDI & PAC |  PBI & pac ; 
 PFJ <= PDJ & PAC |  PBJ & pac ; 
 PBA <= NAA ; 
 PBB <= NAB ; 
 PBC <= NAC ; 
 PBE <= NAE ; 
 PBI <= NAI ; 
 PBM <= NAM ; 
 PCA <= NBA ; 
 PCE <= NBE ; 
 PCI <= NBI ; 
 PCM <= NBM ; 
 PDE <= nae ; 
 PDI <= nai ; 
 PDM <= nam ; 
 PEA <= nba ; 
 PEE <= nbe ; 
 PEI <= nbi ; 
 PEM <= nbm ; 
 GRC <= END ; 
 PAF <=  NED & NXB & NXC & NXD & NXE  |  NHE & NXC & NXD & NXE  |  NIE & NXD & NXE  |  NJE & NXE & NXE  |  NKE  ; 
 PCB <= NBB & nkb |  nbb & NKB ; 
 PCC <= NBC & nkc |  nbc & NKC ; 
 PCD <= NBD & nkd |  nbd & NKD ; 
 PCF <= NBF & nlb |  nbf & NLB ; 
 PCG <= NBG & nlc |  nbg & NLC ; 
 PCH <= NBH & nld |  nbh & NLD ; 
 PEO <= NBO & nvc |  nbo & NVC ; 
 PEN <= NBN & nvb |  nbn & NVB ; 
 PAH <=  NIE & NXD & NXE & NXF & NXG  |  NJE & NXE & NXF & NXG  |  NKE & NXF & NXG  |  NLE & NXG & NXG  |  NME  ; 
 MAF <=  LGA & lgc & lhb  |  lga & LGC & lhb  |  lga & lgc & LHB  |  LGA & LGC & LHB  ;
 mcf <=  LGA & lgc & lhb  |  lga & LGC & lhb  |  lga & lgc & LHB  |  lga & lgc & lhb  ;
 QAA <= IHA ; 
 QAB <= QAA ; 
 QAC <= QAB ; 
 QAD <= QAC ; 
 QAE <= QAD ; 
 QAF <= QAE ; 
 QAG <= QAF ; 
 QAH <= QAG ; 
 MAG <=  LHA & lhc & lib  |  lha & LHC & lib  |  lha & lhc & LIB  |  LHA & LHC & LIB  ;
 mcg <=  LHA & lhc & lib  |  lha & LHC & lib  |  lha & lhc & LIB  |  lha & lhc & lib  ;
 OEA <= IEA ; 
 OEB <= IEB ; 
 OEC <= IEC ; 
 OED <= IED ; 
 OEE <= IEE ; 
 OEF <= IEF ; 
 OFA <= IEA ; 
 OFB <= IEB ; 
 OFC <= IEC ; 
 OFD <= IED ; 
 OFE <= IEE ; 
 OFF <= IEF ; 
 MAH <=  LIA & lic & ljb  |  lia & LIC & ljb  |  lia & lic & LJB  |  LIA & LIC & LJB  ;
 mch <=  LIA & lic & ljb  |  lia & LIC & ljb  |  lia & lic & LJB  |  lia & lic & ljb  ;
 GYB <= EGB & EHA ; 
 ohc <= EGB & iec ; 
 ohd <= EGB & ied ; 
 ohe <= EGB & iee ; 
 oga <= iea ; 
 ogb <= ieb ; 
 ogc <= iec ; 
 ogd <= ied ; 
 oge <= iee ; 
 ogf <= ief ; 
 oha <= iea ; 
 ohb <= ieb ; 
 MAI <=  LJA & ljc & lkb  |  lja & LJC & lkb  |  lja & ljc & LKB  |  LJA & LJC & LKB  ;
 mci <=  LJA & ljc & lkb  |  lja & LJC & lkb  |  lja & ljc & LKB  |  lja & ljc & lkb  ;
 oig <= ifg ; 
 okg <= ifg ; 
 omg <= ifg ; 
 oog <= ifg ; 
 QAI <= QAH ; 
 QAJ <= QAI ; 
 QAK <= QAJ ; 
 NBQ <= MEC ; 
 MAJ <=  LKA & lkc & llb  |  lka & LKC & llb  |  lka & lkc & LLB  |  LKA & LKC & LLB  ;
 mcj <=  LKA & lkc & llb  |  lka & LKC & llb  |  lka & lkc & LLB  |  lka & lkc & llb  ;
 ACE <= AAE ; 
 ACF <= AAF ; 
 ACG <= AAG ; 
 ACH <= AAH ; 
 ACI <= AAI ; 
 ACJ <= AAJ ; 
 ACK <= AAK ; 
 ACL <= AAL ; 
 ACM <= AAM ; 
 ACN <= AAN ; 
 ACO <= AAO ; 
 ACP <= AAP ; 
 MAK <=  LLA & llc & lmb  |  lla & LLC & lmb  |  lla & llc & LMB  |  LLA & LLC & LMB  ;
 mck <=  LLA & llc & lmb  |  lla & LLC & lmb  |  lla & llc & LMB  |  lla & llc & lmb  ;
 PCJ <= NBJ & nmb |  nbj & NMB ; 
 PCK <= NBK & nmc |  nbk & NMC ; 
 PCL <= NBL & nmd |  nbl & NMD ; 
 PCN <= NBN & nnb |  nbn & NNB ; 
 PCO <= NBO & nnc |  nbo & NNC ; 
 PCP <= NBP & nnd |  nbp & NND ; 
 MAL <=  LMA & lmc & lnb  |  lma & LMC & lnb  |  lma & lmc & LNB  |  LMA & LMC & LNB  ;
 mcl <=  LMA & lmc & lnb  |  lma & LMC & lnb  |  lma & lmc & LNB  |  lma & lmc & lnb  ;
 MAM <=  LNA & lnc & lob  |  lna & LNC & lob  |  lna & lnc & LOB  |  LNA & LNC & LOB  ;
 mcm <=  LNA & lnc & lob  |  lna & LNC & lob  |  lna & lnc & LOB  |  lna & lnc & lob  ;
 DRA <=  CAN & cbn & ccm  |  can & CBN & ccm  |  can & cbn & CCM  |  CAN & CBN & CCM  ;
 drb <=  CAN & cbn & ccm  |  can & CBN & ccm  |  can & cbn & CCM  |  can & cbn & ccm  ;
 BAG <= IAG & tee |  BAG & TEE ; 
 BAH <= IAH & tee |  BAH & TEE ; 
 BAO <= IAO & tef |  BAO & TEF ; 
 BAP <= IAP & tef |  BAP & TEF ; 
 BBO <= IBO & teh |  BBO & TEH ; 
 BBP <= IBP & teh |  BBP & TEH ; 
 DRC <=  CDM & cel & cfl  |  cdm & CEL & cfl  |  cdm & cel & CFL  |  CDM & CEL & CFL  ;
 drd <=  CDM & cel & cfl  |  cdm & CEL & cfl  |  cdm & cel & CFL  |  cdm & cel & cfl  ;
 BBG <= IBG & teg |  BBG & TEG ; 
 BBH <= IBH & teg |  BBH & TEG ; 
 KZE <= JZC ; 
 KZF <= JZD ; 
 DRE <=  CGK & chk & cij  |  cgk & CHK & cij  |  cgk & chk & CIJ  |  CGK & CHK & CIJ  ;
 drf <=  CGK & chk & cij  |  cgk & CHK & cij  |  cgk & chk & CIJ  |  cgk & chk & cij  ;
 DRG <=  CJJ & cki & cli  |  cjj & CKI & cli  |  cjj & cki & CLI  |  CJJ & CKI & CLI  ;
 drh <=  CJJ & cki & cli  |  cjj & CKI & cli  |  cjj & cki & CLI  |  cjj & cki & cli  ;
 OJK <= IGD ; 
 OLK <= IGD ; 
 ONK <= IGD ; 
 OPK <= IGD ; 
 DRI <=  CMH & cnh & cog  |  cmh & CNH & cog  |  cmh & cnh & COG  |  CMH & CNH & COG  ;
 drj <=  CMH & cnh & cog  |  cmh & CNH & cog  |  cmh & cnh & COG  |  cmh & cnh & cog  ;
 OJL <= IGE ; 
 OLL <= IGE ; 
 ONL <= IGE ; 
 OPL <= IGE ; 
 OJF <= IFF ; 
 OLF <= IFF ; 
 ONF <= IFF ; 
 OPF <= IFF ; 
 MBM <= LZJ ; 
 DRK <=  CPG & cqf & crf  |  cpg & CQF & crf  |  cpg & cqf & CRF  |  CPG & CQF & CRF  ;
 drl <=  CPG & cqf & crf  |  cpg & CQF & crf  |  cpg & cqf & CRF  |  cpg & cqf & crf  ;
 OJJ <= IGC ; 
 OLJ <= IGC ; 
 ONJ <= IGC ; 
 OPJ <= IGC ; 
 DRM <=  CSE & cte & cud  |  cse & CTE & cud  |  cse & cte & CUD  |  CSE & CTE & CUD  ;
 drn <=  CSE & cte & cud  |  cse & CTE & cud  |  cse & cte & CUD  |  cse & cte & cud  ;
 ACQ <= AAQ ; 
 PGN <=  PCN & pah & pam  |  PEN & PAH  |  PEN & PAM  ; 
 PGP <=  PCP & pah & pam  |  PEP & PAH  |  PEP & PAM  ; 
 DRO <=  CVD & cwc & cxc  |  cvd & CWC & cxc  |  cvd & cwc & CXC  |  CVD & CWC & CXC  ;
 drp <=  CVD & cwc & cxc  |  cvd & CWC & cxc  |  cvd & cwc & CXC  |  cvd & cwc & cxc  ;
 TFA <= QAI ; 
 TFB <= QAI ; 
 TFC <= QAI ; 
 TFD <= QAI ; 
 MEB <= LDB & ldd |  ldb & LDD ; 
 GYA <= EHA & egb |  eha & EGB ; 
 GZA <= EGA & efb |  ega & EFB ; 
 GZB <= EFB & EGA ; 
 GZE <= EEB & EFA ; 
 MDN <= LZO ; 
 PAG <=  NHE & NXC & NXD & NXE & NXF  |  NIE & NXD & NXE & NXF  |  NJE & NXE & NXF  |  NKE & NXF & NXF  |  NLE  ; 
 ADA <= ABA ; 
 ADB <= ABB ; 
 ADC <= ABC ; 
 ADD <= ABD ; 
 ADE <= ABE ; 
 ADF <= ABF ; 
 ADG <= ABG ; 
 ADH <= ABH ; 
 pai <=  nxc  |  nxd  |  nxe  |  nxf  |  nxg  ; 
 ADI <= ABI ; 
 ADJ <= ABJ ; 
 ADK <= ABK ; 
 ADL <= ABL ; 
 PEF <= NBF & ntb |  nbf & NTB ; 
 ADM <= ABM ; 
 ADN <= ABN ; 
 ADO <= ABO ; 
 ADP <= ABP ; 
 ACA <= AAA ; 
 ACB <= AAB ; 
 ACC <= AAC ; 
 ACD <= AAD ; 
 MAA <=  LBA & lbc & lcb  |  lba & LBC & lcb  |  lba & lbc & LCB  |  LBA & LBC & LCB  ;
 mca <=  LBA & lbc & lcb  |  lba & LBC & lcb  |  lba & lbc & LCB  |  lba & lbc & lcb  ;
 PGJ <=  PCJ & pag & pak  |  PEJ & PAG  |  PEJ & PAK  ; 
 PGL <=  PCL & pag & pak  |  PEL & PAG  |  PEL & PAK  ; 
 OJM <= IGF ; 
 OLM <= IGF ; 
 ONM <= IGF ; 
 OPM <= IGF ; 
 end 
end module
