module fa( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFF, 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 IHM, 
 IHN, 
 IHO, 
 IHP, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IKA, 
 ILA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OAR, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OIA, 
 OJA, 
 OJB, 
 OJC, 
OKA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFF; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 input IHM; 
 input IHN; 
 input IHO; 
 input IHP; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IKA; 
 input ILA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OAR; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OIA; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OKA; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  aea ;
reg  aeb ;
reg  aec ;
reg  aed ;
reg  aee ;
reg  aef ;
reg  aeg ;
reg  aeh ;
reg  aei ;
reg  aej ;
reg  aek ;
reg  ael ;
reg  aem ;
reg  aen ;
reg  aeo ;
reg  aep ;
reg  afa ;
reg  afb ;
reg  afc ;
reg  afd ;
reg  afe ;
reg  aff ;
reg  afg ;
reg  afh ;
reg  afi ;
reg  afj ;
reg  afk ;
reg  afl ;
reg  afm ;
reg  afn ;
reg  afo ;
reg  afp ;
reg  aga ;
reg  agb ;
reg  agc ;
reg  agd ;
reg  age ;
reg  agf ;
reg  agg ;
reg  agh ;
reg  agi ;
reg  agj ;
reg  agk ;
reg  agl ;
reg  agm ;
reg  agn ;
reg  ago ;
reg  agp ;
reg  aha ;
reg  ahb ;
reg  ahc ;
reg  ahd ;
reg  ahe ;
reg  ahf ;
reg  ahg ;
reg  ahh ;
reg  ahi ;
reg  ahj ;
reg  ahk ;
reg  ahl ;
reg  ahm ;
reg  ahn ;
reg  aho ;
reg  ahp ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  caa ;
reg  cab ;
reg  cac ;
reg  cad ;
reg  cae ;
reg  caf ;
reg  cag ;
reg  cah ;
reg  cai ;
reg  caj ;
reg  cak ;
reg  cal ;
reg  cam ;
reg  can ;
reg  cao ;
reg  cba ;
reg  cbb ;
reg  cbc ;
reg  cbg ;
reg  cbh ;
reg  DCB ;
reg  DCC ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FBA ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FBE ;
reg  FBF ;
reg  FBG ;
reg  FBH ;
reg  FBI ;
reg  FBJ ;
reg  FBK ;
reg  FBL ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FIE ;
reg  FIF ;
reg  FIG ;
reg  FIH ;
reg  FII ;
reg  FIJ ;
reg  FIK ;
reg  FIL ;
reg  FIM ;
reg  FIN ;
reg  FIO ;
reg  FIP ;
reg  FJA ;
reg  FJB ;
reg  FJC ;
reg  FJD ;
reg  FJE ;
reg  FJF ;
reg  FJG ;
reg  FJH ;
reg  FJI ;
reg  FJJ ;
reg  FJK ;
reg  FJL ;
reg  FJM ;
reg  FJN ;
reg  FJO ;
reg  FJP ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FKE ;
reg  FKF ;
reg  FKG ;
reg  FKH ;
reg  FKI ;
reg  FKJ ;
reg  FKK ;
reg  FKL ;
reg  FKM ;
reg  FKN ;
reg  FKO ;
reg  FKP ;
reg  FLA ;
reg  FLB ;
reg  FLC ;
reg  FLD ;
reg  FLE ;
reg  FLF ;
reg  FLG ;
reg  FLH ;
reg  FLI ;
reg  FLJ ;
reg  FLK ;
reg  FLL ;
reg  FLM ;
reg  FLN ;
reg  FLO ;
reg  FLP ;
reg  FMA ;
reg  FMB ;
reg  FMC ;
reg  FMD ;
reg  FME ;
reg  FMF ;
reg  FMG ;
reg  FMH ;
reg  FMI ;
reg  FMJ ;
reg  FMK ;
reg  FML ;
reg  FMM ;
reg  FMN ;
reg  FMO ;
reg  FMP ;
reg  FNA ;
reg  FNB ;
reg  FNC ;
reg  FND ;
reg  FNE ;
reg  FNF ;
reg  FNG ;
reg  FNH ;
reg  FNI ;
reg  FNJ ;
reg  FNK ;
reg  FNL ;
reg  FNM ;
reg  FNN ;
reg  FNO ;
reg  FNP ;
reg  FOA ;
reg  FOB ;
reg  FOC ;
reg  FOD ;
reg  FOE ;
reg  FOF ;
reg  FOG ;
reg  FOH ;
reg  FOI ;
reg  FOJ ;
reg  FOK ;
reg  FOL ;
reg  FOM ;
reg  FON ;
reg  FOO ;
reg  FOP ;
reg  FPA ;
reg  FPB ;
reg  FPC ;
reg  FPD ;
reg  FPE ;
reg  FPF ;
reg  FPG ;
reg  FPH ;
reg  FPI ;
reg  FPJ ;
reg  FPK ;
reg  FPL ;
reg  FPM ;
reg  FPN ;
reg  FPO ;
reg  FPP ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GAI ;
reg  GAJ ;
reg  GAK ;
reg  GAL ;
reg  GAM ;
reg  GAN ;
reg  GAO ;
reg  gap ;
reg  gaq ;
reg  gba ;
reg  gca ;
reg  HBK ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  KAQ ;
reg  kar ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KBI ;
reg  KBJ ;
reg  KBK ;
reg  KBL ;
reg  KBM ;
reg  KBN ;
reg  KBO ;
reg  KBP ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  KCD ;
reg  KCE ;
reg  KCF ;
reg  KCG ;
reg  KCH ;
reg  KCI ;
reg  KCJ ;
reg  KCK ;
reg  KCL ;
reg  KCM ;
reg  KCN ;
reg  KCO ;
reg  KCP ;
reg  kda ;
reg  kdb ;
reg  kdc ;
reg  kdd ;
reg  kde ;
reg  kdf ;
reg  kdg ;
reg  kdh ;
reg  kdi ;
reg  kdj ;
reg  kdk ;
reg  kdl ;
reg  kdm ;
reg  kdn ;
reg  kdo ;
reg  kdp ;
reg  kea ;
reg  keb ;
reg  kec ;
reg  ked ;
reg  kee ;
reg  kef ;
reg  keg ;
reg  keh ;
reg  kei ;
reg  kej ;
reg  kek ;
reg  kel ;
reg  kem ;
reg  ken ;
reg  keo ;
reg  kep ;
reg  kfa ;
reg  kfb ;
reg  kfc ;
reg  kfd ;
reg  kfe ;
reg  kff ;
reg  kfg ;
reg  kfh ;
reg  kfi ;
reg  kfj ;
reg  kfk ;
reg  kfl ;
reg  kfm ;
reg  kfn ;
reg  kfo ;
reg  kfp ;
reg  kja ;
reg  kjb ;
reg  kjc ;
reg  kjd ;
reg  kje ;
reg  kjf ;
reg  kjg ;
reg  kjh ;
reg  kji ;
reg  kjj ;
reg  kjk ;
reg  kjl ;
reg  kjm ;
reg  kjn ;
reg  kjo ;
reg  kjp ;
reg  kka ;
reg  kkb ;
reg  kkc ;
reg  kkd ;
reg  kke ;
reg  kkf ;
reg  kkg ;
reg  kkh ;
reg  kki ;
reg  kkj ;
reg  kkk ;
reg  kkl ;
reg  kkm ;
reg  kkn ;
reg  kko ;
reg  kkp ;
reg  KLD ;
reg  KLH ;
reg  KLI ;
reg  KLJ ;
reg  KLK ;
reg  KLL ;
reg  KLM ;
reg  KLN ;
reg  KLO ;
reg  KLP ;
reg  KMA ;
reg  KMB ;
reg  KMC ;
reg  KMD ;
reg  KME ;
reg  KMF ;
reg  KMG ;
reg  KMH ;
reg  KMI ;
reg  KMJ ;
reg  KMK ;
reg  KML ;
reg  KMM ;
reg  KMN ;
reg  KMO ;
reg  KMP ;
reg  KNA ;
reg  KNB ;
reg  KNC ;
reg  KND ;
reg  KNE ;
reg  KNI ;
reg  KNJ ;
reg  KNK ;
reg  KNL ;
reg  KNM ;
reg  KOA ;
reg  KOB ;
reg  KOC ;
reg  KOD ;
reg  KOE ;
reg  KOF ;
reg  KOG ;
reg  KOH ;
reg  KOI ;
reg  KOJ ;
reg  KOK ;
reg  KOL ;
reg  KOM ;
reg  KON ;
reg  KOO ;
reg  KOP ;
reg  KPA ;
reg  KPB ;
reg  KPC ;
reg  KPD ;
reg  KPE ;
reg  KPI ;
reg  KPJ ;
reg  KPK ;
reg  KPL ;
reg  KPM ;
reg  KQL ;
reg  KQM ;
reg  oaa ;
reg  oab ;
reg  oac ;
reg  oad ;
reg  oae ;
reg  oaf ;
reg  oag ;
reg  oah ;
reg  oai ;
reg  oaj ;
reg  oak ;
reg  oal ;
reg  oam ;
reg  oan ;
reg  oao ;
reg  oap ;
reg  oar ;
reg  oba ;
reg  obb ;
reg  obc ;
reg  obd ;
reg  obe ;
reg  obf ;
reg  obg ;
reg  obh ;
reg  obi ;
reg  obj ;
reg  obk ;
reg  obl ;
reg  obm ;
reg  obn ;
reg  obo ;
reg  obp ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  odk ;
reg  odl ;
reg  odm ;
reg  odn ;
reg  odo ;
reg  odp ;
reg  oea ;
reg  oeb ;
reg  oec ;
reg  oed ;
reg  oee ;
reg  oef ;
reg  oeg ;
reg  oeh ;
reg  oei ;
reg  oej ;
reg  oek ;
reg  oel ;
reg  oem ;
reg  oen ;
reg  oeo ;
reg  oep ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  ofe ;
reg  off ;
reg  ofg ;
reg  ofh ;
reg  ofi ;
reg  ofj ;
reg  ofk ;
reg  ofl ;
reg  ofm ;
reg  ofn ;
reg  ofo ;
reg  ofp ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OHA ;
reg  OIA ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  oka ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  qae ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  qbf ;
reg  qbg ;
reg  qbh ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  QCE ;
reg  QCF ;
reg  QCG ;
reg  QCH ;
reg  QCI ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QDF ;
reg  QDG ;
reg  QDH ;
reg  qdi ;
reg  qdj ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  QED ;
reg  QEE ;
reg  QEF ;
reg  QEG ;
reg  QEH ;
reg  QEI ;
reg  QEJ ;
reg  QEK ;
reg  qfa ;
reg  qfb ;
reg  qfc ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  QGE ;
reg  QGF ;
reg  qgg ;
reg  qgh ;
reg  qgi ;
reg  qgj ;
reg  QHA ;
reg  QHB ;
reg  QHC ;
reg  QIA ;
reg  QIB ;
reg  qja ;
reg  QJM ;
reg  qka ;
reg  qkb ;
reg  QKC ;
reg  qkd ;
reg  qke ;
reg  qkf ;
reg  qkg ;
reg  qkh ;
reg  qki ;
reg  qkj ;
reg  qkk ;
reg  qkl ;
reg  qxa ;
reg  qxb ;
reg  qxc ;
reg  qxd ;
reg  qxe ;
reg  qxf ;
reg  qxg ;
reg  qxh ;
reg  qxi ;
reg  QXJ ;
reg  QXK ;
reg  QXL ;
reg  qxm ;
reg  QYA ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  RAI ;
reg  RAJ ;
reg  RAK ;
reg  RAL ;
reg  RAM ;
reg  RAN ;
reg  RAO ;
reg  RAP ;
reg  RBA ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  RBH ;
reg  RBI ;
reg  RBJ ;
reg  RBK ;
reg  RBL ;
reg  RBM ;
reg  RBN ;
reg  RBO ;
reg  RBP ;
reg  RCA ;
reg  RCB ;
reg  RCC ;
reg  RCD ;
reg  RCE ;
reg  RCF ;
reg  RCG ;
reg  RCH ;
reg  RCI ;
reg  RCJ ;
reg  RCK ;
reg  RCL ;
reg  RCM ;
reg  RCN ;
reg  RCO ;
reg  RCP ;
reg  taa ;
reg  tab ;
reg  tac ;
reg  tad ;
reg  tba ;
reg  tca ;
reg  tcb ;
reg  tcc ;
reg  tcd ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TEA ;
reg  TFA ;
reg  TFB ;
reg  tga ;
reg  tgb ;
reg  tgc ;
reg  tgd ;
reg  tge ;
reg  tgf ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TMD ;
reg  TME ;
reg  TMF ;
reg  TNA ;
reg  TNB ;
reg  TNC ;
reg  TND ;
reg  TNE ;
reg  TNF ;
reg  TOA ;
reg  TOB ;
reg  TOC ;
reg  TOD ;
reg  TOE ;
reg  TOF ;
reg  TPA ;
reg  TPB ;
reg  TPC ;
reg  TPD ;
reg  TPE ;
reg  TPF ;
reg  TQA ;
reg  TQB ;
reg  TQC ;
reg  TQD ;
reg  TQE ;
reg  TQF ;
reg  TQG ;
reg  TQH ;
reg  TQI ;
reg  TQJ ;
reg  TQK ;
reg  TQL ;
reg  tqm ;
reg  tqn ;
reg  tqo ;
reg  TRA ;
reg  TRB ;
reg  TRC ;
reg  TRD ;
reg  TRE ;
reg  TRF ;
reg  TRG ;
reg  TRH ;
reg  TRI ;
reg  TRJ ;
reg  TRK ;
reg  TRL ;
reg  TSA ;
reg  TSB ;
reg  TSC ;
reg  TSD ;
reg  TSE ;
reg  TSF ;
reg  TSG ;
reg  TSH ;
reg  TSI ;
reg  TSJ ;
reg  TSK ;
reg  TSL ;
reg  TTA ;
reg  TTB ;
reg  TTC ;
reg  TTD ;
reg  TTE ;
reg  TTF ;
reg  TTG ;
reg  TTH ;
reg  TTI ;
reg  TTJ ;
reg  TTK ;
reg  TTL ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  AEA ;
wire  AEB ;
wire  AEC ;
wire  AED ;
wire  AEE ;
wire  AEF ;
wire  AEG ;
wire  AEH ;
wire  AEI ;
wire  AEJ ;
wire  AEK ;
wire  AEL ;
wire  AEM ;
wire  AEN ;
wire  AEO ;
wire  AEP ;
wire  AFA ;
wire  AFB ;
wire  AFC ;
wire  AFD ;
wire  AFE ;
wire  AFF ;
wire  AFG ;
wire  AFH ;
wire  AFI ;
wire  AFJ ;
wire  AFK ;
wire  AFL ;
wire  AFM ;
wire  AFN ;
wire  AFO ;
wire  AFP ;
wire  AGA ;
wire  AGB ;
wire  AGC ;
wire  AGD ;
wire  AGE ;
wire  AGF ;
wire  AGG ;
wire  AGH ;
wire  AGI ;
wire  AGJ ;
wire  AGK ;
wire  AGL ;
wire  AGM ;
wire  AGN ;
wire  AGO ;
wire  AGP ;
wire  AHA ;
wire  AHB ;
wire  AHC ;
wire  AHD ;
wire  AHE ;
wire  AHF ;
wire  AHG ;
wire  AHH ;
wire  AHI ;
wire  AHJ ;
wire  AHK ;
wire  AHL ;
wire  AHM ;
wire  AHN ;
wire  AHO ;
wire  AHP ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  CAA ;
wire  CAB ;
wire  CAC ;
wire  CAD ;
wire  CAE ;
wire  CAF ;
wire  CAG ;
wire  CAH ;
wire  CAI ;
wire  CAJ ;
wire  CAK ;
wire  CAL ;
wire  CAM ;
wire  CAN ;
wire  CAO ;
wire  CBA ;
wire  CBB ;
wire  CBC ;
wire  CBG ;
wire  CBH ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  dae ;
wire  DAE ;
wire  daf ;
wire  DAF ;
wire  dag ;
wire  DAG ;
wire  dah ;
wire  DAH ;
wire  dai ;
wire  DAI ;
wire  daj ;
wire  DAJ ;
wire  dak ;
wire  DAK ;
wire  dal ;
wire  DAL ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dbe ;
wire  DBE ;
wire  dbf ;
wire  DBF ;
wire  dbg ;
wire  DBG ;
wire  dbh ;
wire  DBH ;
wire  dbi ;
wire  DBI ;
wire  dbj ;
wire  DBJ ;
wire  dbk ;
wire  DBK ;
wire  dbl ;
wire  DBL ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  DCD ;
wire  dce ;
wire  DCE ;
wire  dcf ;
wire  DCF ;
wire  ddg ;
wire  DDG ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fba ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fbe ;
wire  fbf ;
wire  fbg ;
wire  fbh ;
wire  fbi ;
wire  fbj ;
wire  fbk ;
wire  fbl ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fie ;
wire  fif ;
wire  fig ;
wire  fih ;
wire  fii ;
wire  fij ;
wire  fik ;
wire  fil ;
wire  fim ;
wire  fin ;
wire  fio ;
wire  fip ;
wire  fja ;
wire  fjb ;
wire  fjc ;
wire  fjd ;
wire  fje ;
wire  fjf ;
wire  fjg ;
wire  fjh ;
wire  fji ;
wire  fjj ;
wire  fjk ;
wire  fjl ;
wire  fjm ;
wire  fjn ;
wire  fjo ;
wire  fjp ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fke ;
wire  fkf ;
wire  fkg ;
wire  fkh ;
wire  fki ;
wire  fkj ;
wire  fkk ;
wire  fkl ;
wire  fkm ;
wire  fkn ;
wire  fko ;
wire  fkp ;
wire  fla ;
wire  flb ;
wire  flc ;
wire  fld ;
wire  fle ;
wire  flf ;
wire  flg ;
wire  flh ;
wire  fli ;
wire  flj ;
wire  flk ;
wire  fll ;
wire  flm ;
wire  fln ;
wire  flo ;
wire  flp ;
wire  fma ;
wire  fmb ;
wire  fmc ;
wire  fmd ;
wire  fme ;
wire  fmf ;
wire  fmg ;
wire  fmh ;
wire  fmi ;
wire  fmj ;
wire  fmk ;
wire  fml ;
wire  fmm ;
wire  fmn ;
wire  fmo ;
wire  fmp ;
wire  fna ;
wire  fnb ;
wire  fnc ;
wire  fnd ;
wire  fne ;
wire  fnf ;
wire  fng ;
wire  fnh ;
wire  fni ;
wire  fnj ;
wire  fnk ;
wire  fnl ;
wire  fnm ;
wire  fnn ;
wire  fno ;
wire  fnp ;
wire  foa ;
wire  fob ;
wire  foc ;
wire  fod ;
wire  foe ;
wire  fof ;
wire  fog ;
wire  foh ;
wire  foi ;
wire  foj ;
wire  fok ;
wire  fol ;
wire  fom ;
wire  fon ;
wire  foo ;
wire  fop ;
wire  fpa ;
wire  fpb ;
wire  fpc ;
wire  fpd ;
wire  fpe ;
wire  fpf ;
wire  fpg ;
wire  fph ;
wire  fpi ;
wire  fpj ;
wire  fpk ;
wire  fpl ;
wire  fpm ;
wire  fpn ;
wire  fpo ;
wire  fpp ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gai ;
wire  gaj ;
wire  gak ;
wire  gal ;
wire  gam ;
wire  gan ;
wire  gao ;
wire  GAP ;
wire  GAQ ;
wire  GBA ;
wire  GCA ;
wire  haa ;
wire  HAA ;
wire  hab ;
wire  HAB ;
wire  hac ;
wire  HAC ;
wire  had ;
wire  HAD ;
wire  hae ;
wire  HAE ;
wire  haf ;
wire  HAF ;
wire  hag ;
wire  HAG ;
wire  hah ;
wire  HAH ;
wire  hai ;
wire  HAI ;
wire  haj ;
wire  HAJ ;
wire  hak ;
wire  HAK ;
wire  hal ;
wire  HAL ;
wire  ham ;
wire  HAM ;
wire  han ;
wire  HAN ;
wire  hao ;
wire  HAO ;
wire  hap ;
wire  HAP ;
wire  hba ;
wire  HBA ;
wire  hbb ;
wire  HBB ;
wire  hbc ;
wire  HBC ;
wire  hbd ;
wire  HBD ;
wire  hbe ;
wire  HBE ;
wire  hbf ;
wire  HBF ;
wire  hbg ;
wire  HBG ;
wire  hbh ;
wire  HBH ;
wire  hbi ;
wire  HBI ;
wire  hbj ;
wire  HBJ ;
wire  hbk ;
wire  hbl ;
wire  HBL ;
wire  hbm ;
wire  HBM ;
wire  hbn ;
wire  HBN ;
wire  hbo ;
wire  HBO ;
wire  hbp ;
wire  HBP ;
wire  hca ;
wire  HCA ;
wire  hcb ;
wire  HCB ;
wire  hcc ;
wire  HCC ;
wire  hcd ;
wire  HCD ;
wire  hce ;
wire  HCE ;
wire  hcf ;
wire  HCF ;
wire  hcg ;
wire  HCG ;
wire  hch ;
wire  HCH ;
wire  hci ;
wire  HCI ;
wire  hcj ;
wire  HCJ ;
wire  hck ;
wire  HCK ;
wire  hcl ;
wire  HCL ;
wire  hcm ;
wire  HCM ;
wire  hcn ;
wire  HCN ;
wire  hco ;
wire  HCO ;
wire  hcp ;
wire  HCP ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iff ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  ihm ;
wire  ihn ;
wire  iho ;
wire  ihp ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ika ;
wire  ila ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jca ;
wire  JCA ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jfc ;
wire  JFC ;
wire  jgc ;
wire  JGC ;
wire  jhc ;
wire  JHC ;
wire  jia ;
wire  JIA ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  kaq ;
wire  KAR ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kbi ;
wire  kbj ;
wire  kbk ;
wire  kbl ;
wire  kbm ;
wire  kbn ;
wire  kbo ;
wire  kbp ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  kcd ;
wire  kce ;
wire  kcf ;
wire  kcg ;
wire  kch ;
wire  kci ;
wire  kcj ;
wire  kck ;
wire  kcl ;
wire  kcm ;
wire  kcn ;
wire  kco ;
wire  kcp ;
wire  KDA ;
wire  KDB ;
wire  KDC ;
wire  KDD ;
wire  KDE ;
wire  KDF ;
wire  KDG ;
wire  KDH ;
wire  KDI ;
wire  KDJ ;
wire  KDK ;
wire  KDL ;
wire  KDM ;
wire  KDN ;
wire  KDO ;
wire  KDP ;
wire  KEA ;
wire  KEB ;
wire  KEC ;
wire  KED ;
wire  KEE ;
wire  KEF ;
wire  KEG ;
wire  KEH ;
wire  KEI ;
wire  KEJ ;
wire  KEK ;
wire  KEL ;
wire  KEM ;
wire  KEN ;
wire  KEO ;
wire  KEP ;
wire  KFA ;
wire  KFB ;
wire  KFC ;
wire  KFD ;
wire  KFE ;
wire  KFF ;
wire  KFG ;
wire  KFH ;
wire  KFI ;
wire  KFJ ;
wire  KFK ;
wire  KFL ;
wire  KFM ;
wire  KFN ;
wire  KFO ;
wire  KFP ;
wire  KJA ;
wire  KJB ;
wire  KJC ;
wire  KJD ;
wire  KJE ;
wire  KJF ;
wire  KJG ;
wire  KJH ;
wire  KJI ;
wire  KJJ ;
wire  KJK ;
wire  KJL ;
wire  KJM ;
wire  KJN ;
wire  KJO ;
wire  KJP ;
wire  KKA ;
wire  KKB ;
wire  KKC ;
wire  KKD ;
wire  KKE ;
wire  KKF ;
wire  KKG ;
wire  KKH ;
wire  KKI ;
wire  KKJ ;
wire  KKK ;
wire  KKL ;
wire  KKM ;
wire  KKN ;
wire  KKO ;
wire  KKP ;
wire  kld ;
wire  klh ;
wire  kli ;
wire  klj ;
wire  klk ;
wire  kll ;
wire  klm ;
wire  kln ;
wire  klo ;
wire  klp ;
wire  kma ;
wire  kmb ;
wire  kmc ;
wire  kmd ;
wire  kme ;
wire  kmf ;
wire  kmg ;
wire  kmh ;
wire  kmi ;
wire  kmj ;
wire  kmk ;
wire  kml ;
wire  kmm ;
wire  kmn ;
wire  kmo ;
wire  kmp ;
wire  kna ;
wire  knb ;
wire  knc ;
wire  knd ;
wire  kne ;
wire  kni ;
wire  knj ;
wire  knk ;
wire  knl ;
wire  knm ;
wire  koa ;
wire  kob ;
wire  koc ;
wire  kod ;
wire  koe ;
wire  kof ;
wire  kog ;
wire  koh ;
wire  koi ;
wire  koj ;
wire  kok ;
wire  kol ;
wire  kom ;
wire  kon ;
wire  koo ;
wire  kop ;
wire  kpa ;
wire  kpb ;
wire  kpc ;
wire  kpd ;
wire  kpe ;
wire  kpi ;
wire  kpj ;
wire  kpk ;
wire  kpl ;
wire  kpm ;
wire  kql ;
wire  kqm ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lac ;
wire  LAC ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  LAE ;
wire  laf ;
wire  LAF ;
wire  lag ;
wire  LAG ;
wire  lah ;
wire  LAH ;
wire  lai ;
wire  LAI ;
wire  laj ;
wire  LAJ ;
wire  lak ;
wire  LAK ;
wire  lal ;
wire  LAL ;
wire  lam ;
wire  LAM ;
wire  lan ;
wire  LAN ;
wire  lao ;
wire  LAO ;
wire  lap ;
wire  LAP ;
wire  lar ;
wire  LAR ;
wire  lba ;
wire  LBA ;
wire  lbb ;
wire  LBB ;
wire  lbc ;
wire  LBC ;
wire  lbd ;
wire  LBD ;
wire  lbe ;
wire  LBE ;
wire  lbf ;
wire  LBF ;
wire  lbg ;
wire  LBG ;
wire  lbh ;
wire  LBH ;
wire  lbi ;
wire  LBI ;
wire  lbj ;
wire  LBJ ;
wire  lbk ;
wire  LBK ;
wire  lbl ;
wire  LBL ;
wire  lbm ;
wire  LBM ;
wire  lbn ;
wire  LBN ;
wire  lbo ;
wire  LBO ;
wire  lbp ;
wire  LBP ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lcc ;
wire  LCC ;
wire  lcd ;
wire  LCD ;
wire  lce ;
wire  LCE ;
wire  lcf ;
wire  LCF ;
wire  lcg ;
wire  LCG ;
wire  lch ;
wire  LCH ;
wire  lci ;
wire  LCI ;
wire  lcj ;
wire  LCJ ;
wire  lck ;
wire  LCK ;
wire  lcl ;
wire  LCL ;
wire  lcm ;
wire  LCM ;
wire  lcn ;
wire  LCN ;
wire  lco ;
wire  LCO ;
wire  lcp ;
wire  LCP ;
wire  ldc ;
wire  LDC ;
wire  ldd ;
wire  LDD ;
wire  ldh ;
wire  LDH ;
wire  ldi ;
wire  LDI ;
wire  ldj ;
wire  LDJ ;
wire  ldk ;
wire  LDK ;
wire  ldl ;
wire  LDL ;
wire  ldo ;
wire  LDO ;
wire  ldp ;
wire  LDP ;
wire  lea ;
wire  LEA ;
wire  leb ;
wire  LEB ;
wire  lec ;
wire  LEC ;
wire  led ;
wire  LED ;
wire  leh ;
wire  LEH ;
wire  lei ;
wire  LEI ;
wire  lej ;
wire  LEJ ;
wire  lek ;
wire  LEK ;
wire  lel ;
wire  LEL ;
wire  lep ;
wire  LEP ;
wire  lfa ;
wire  LFA ;
wire  lfb ;
wire  LFB ;
wire  lfc ;
wire  LFC ;
wire  lfd ;
wire  LFD ;
wire  lfh ;
wire  LFH ;
wire  lfi ;
wire  LFI ;
wire  lfj ;
wire  LFJ ;
wire  lfk ;
wire  LFK ;
wire  lfl ;
wire  LFL ;
wire  lfp ;
wire  LFP ;
wire  lgi ;
wire  LGI ;
wire  lha ;
wire  LHA ;
wire  lht ;
wire  LHT ;
wire  lia ;
wire  LIA ;
wire  lii ;
wire  LII ;
wire  nba ;
wire  NBA ;
wire  nbb ;
wire  NBB ;
wire  nbc ;
wire  NBC ;
wire  nbd ;
wire  NBD ;
wire  nbe ;
wire  NBE ;
wire  nbf ;
wire  NBF ;
wire  nca ;
wire  NCA ;
wire  ncb ;
wire  NCB ;
wire  ncc ;
wire  NCC ;
wire  OAA ;
wire  OAB ;
wire  OAC ;
wire  OAD ;
wire  OAE ;
wire  OAF ;
wire  OAG ;
wire  OAH ;
wire  OAI ;
wire  OAJ ;
wire  OAK ;
wire  OAL ;
wire  OAM ;
wire  OAN ;
wire  OAO ;
wire  OAP ;
wire  OAR ;
wire  OBA ;
wire  OBB ;
wire  OBC ;
wire  OBD ;
wire  OBE ;
wire  OBF ;
wire  OBG ;
wire  OBH ;
wire  OBI ;
wire  OBJ ;
wire  OBK ;
wire  OBL ;
wire  OBM ;
wire  OBN ;
wire  OBO ;
wire  OBP ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  ODK ;
wire  ODL ;
wire  ODM ;
wire  ODN ;
wire  ODO ;
wire  ODP ;
wire  OEA ;
wire  OEB ;
wire  OEC ;
wire  OED ;
wire  OEE ;
wire  OEF ;
wire  OEG ;
wire  OEH ;
wire  OEI ;
wire  OEJ ;
wire  OEK ;
wire  OEL ;
wire  OEM ;
wire  OEN ;
wire  OEO ;
wire  OEP ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OFE ;
wire  OFF ;
wire  OFG ;
wire  OFH ;
wire  OFI ;
wire  OFJ ;
wire  OFK ;
wire  OFL ;
wire  OFM ;
wire  OFN ;
wire  OFO ;
wire  OFP ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  oha ;
wire  oia ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  OKA ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  QAE ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  QBF ;
wire  QBG ;
wire  QBH ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  qce ;
wire  qcf ;
wire  qcg ;
wire  qch ;
wire  qci ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qdf ;
wire  qdg ;
wire  qdh ;
wire  QDI ;
wire  QDJ ;
wire  qea ;
wire  qeb ;
wire  qec ;
wire  qed ;
wire  qee ;
wire  qef ;
wire  qeg ;
wire  qeh ;
wire  qei ;
wire  qej ;
wire  qek ;
wire  QFA ;
wire  QFB ;
wire  QFC ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  qge ;
wire  qgf ;
wire  QGG ;
wire  QGH ;
wire  QGI ;
wire  QGJ ;
wire  qha ;
wire  qhb ;
wire  qhc ;
wire  qia ;
wire  qib ;
wire  QJA ;
wire  qjm ;
wire  QKA ;
wire  QKB ;
wire  qkc ;
wire  QKD ;
wire  QKE ;
wire  QKF ;
wire  QKG ;
wire  QKH ;
wire  QKI ;
wire  QKJ ;
wire  QKK ;
wire  QKL ;
wire  QXA ;
wire  QXB ;
wire  QXC ;
wire  QXD ;
wire  QXE ;
wire  QXF ;
wire  QXG ;
wire  QXH ;
wire  QXI ;
wire  qxj ;
wire  qxk ;
wire  qxl ;
wire  QXM ;
wire  qya ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  rai ;
wire  raj ;
wire  rak ;
wire  ral ;
wire  ram ;
wire  ran ;
wire  rao ;
wire  rap ;
wire  rba ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  rbh ;
wire  rbi ;
wire  rbj ;
wire  rbk ;
wire  rbl ;
wire  rbm ;
wire  rbn ;
wire  rbo ;
wire  rbp ;
wire  rca ;
wire  rcb ;
wire  rcc ;
wire  rcd ;
wire  rce ;
wire  rcf ;
wire  rcg ;
wire  rch ;
wire  rci ;
wire  rcj ;
wire  rck ;
wire  rcl ;
wire  rcm ;
wire  rcn ;
wire  rco ;
wire  rcp ;
wire  TAA ;
wire  TAB ;
wire  TAC ;
wire  TAD ;
wire  TBA ;
wire  TCA ;
wire  TCB ;
wire  TCC ;
wire  TCD ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tea ;
wire  tfa ;
wire  tfb ;
wire  TGA ;
wire  TGB ;
wire  TGC ;
wire  TGD ;
wire  TGE ;
wire  TGF ;
wire  tha ;
wire  THA ;
wire  thb ;
wire  THB ;
wire  thc ;
wire  THC ;
wire  thd ;
wire  THD ;
wire  the ;
wire  THE ;
wire  thf ;
wire  THF ;
wire  thg ;
wire  THG ;
wire  thh ;
wire  THH ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tmd ;
wire  tme ;
wire  tmf ;
wire  tna ;
wire  tnb ;
wire  tnc ;
wire  tnd ;
wire  tne ;
wire  tnf ;
wire  toa ;
wire  tob ;
wire  toc ;
wire  tod ;
wire  toe ;
wire  tof ;
wire  tpa ;
wire  tpb ;
wire  tpc ;
wire  tpd ;
wire  tpe ;
wire  tpf ;
wire  tqa ;
wire  tqb ;
wire  tqc ;
wire  tqd ;
wire  tqe ;
wire  tqf ;
wire  tqg ;
wire  tqh ;
wire  tqi ;
wire  tqj ;
wire  tqk ;
wire  tql ;
wire  TQM ;
wire  TQN ;
wire  TQO ;
wire  tra ;
wire  trb ;
wire  trc ;
wire  trd ;
wire  tre ;
wire  trf ;
wire  trg ;
wire  trh ;
wire  tri ;
wire  trj ;
wire  trk ;
wire  trl ;
wire  tsa ;
wire  tsb ;
wire  tsc ;
wire  tsd ;
wire  tse ;
wire  tsf ;
wire  tsg ;
wire  tsh ;
wire  tsi ;
wire  tsj ;
wire  tsk ;
wire  tsl ;
wire  tta ;
wire  ttb ;
wire  ttc ;
wire  ttd ;
wire  tte ;
wire  ttf ;
wire  ttg ;
wire  tth ;
wire  tti ;
wire  ttj ;
wire  ttk ;
wire  ttl ;
wire  tua ;
wire  TUA ;
wire  tub ;
wire  TUB ;
wire  tuc ;
wire  TUC ;
wire  tud ;
wire  TUD ;
wire  tue ;
wire  TUE ;
wire  tuf ;
wire  TUF ;
wire  tug ;
wire  TUG ;
wire  tuh ;
wire  TUH ;
wire  tui ;
wire  TUI ;
wire  tuj ;
wire  TUJ ;
wire  tuk ;
wire  TUK ;
wire  tul ;
wire  TUL ;
wire  tva ;
wire  TVA ;
wire  tvb ;
wire  TVB ;
wire  tvc ;
wire  TVC ;
wire  tvd ;
wire  TVD ;
wire  tve ;
wire  TVE ;
wire  tvf ;
wire  TVF ;
wire  tvg ;
wire  TVG ;
wire  tvh ;
wire  TVH ;
wire  tvi ;
wire  TVI ;
wire  tvj ;
wire  TVJ ;
wire  tvk ;
wire  TVK ;
wire  tvl ;
wire  TVL ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign rbi = ~RBI;  //complement 
assign rbj = ~RBJ;  //complement 
assign rbk = ~RBK;  //complement 
assign rbl = ~RBL;  //complement 
assign rci = ~RCI;  //complement 
assign rcj = ~RCJ;  //complement 
assign rck = ~RCK;  //complement 
assign rcl = ~RCL;  //complement 
assign rai = ~RAI;  //complement 
assign raj = ~RAJ;  //complement 
assign fli = ~FLI;  //complement 
assign flj = ~FLJ;  //complement 
assign flk = ~FLK;  //complement 
assign fll = ~FLL;  //complement 
assign rao = ~RAO;  //complement 
assign rap = ~RAP;  //complement 
assign rak = ~RAK;  //complement 
assign ral = ~RAL;  //complement 
assign fpi = ~FPI;  //complement 
assign fpj = ~FPJ;  //complement 
assign fpk = ~FPK;  //complement 
assign fpl = ~FPL;  //complement 
assign KKI = ~kki;  //complement 
assign KKJ = ~kkj;  //complement 
assign KKK = ~kkk;  //complement 
assign KKL = ~kkl;  //complement 
assign KKM = ~kkm;  //complement 
assign KKN = ~kkn;  //complement 
assign KKO = ~kko;  //complement 
assign KKP = ~kkp;  //complement 
assign jeb =  qek & qeg  ; 
assign JEB = ~jeb;  //complement 
assign KJM = ~kjm;  //complement 
assign KJN = ~kjn;  //complement 
assign KJO = ~kjo;  //complement 
assign KJP = ~kjp;  //complement 
assign ram = ~RAM;  //complement 
assign ran = ~RAN;  //complement 
assign fpm = ~FPM;  //complement 
assign fpn = ~FPN;  //complement 
assign fpo = ~FPO;  //complement 
assign fpp = ~FPP;  //complement 
assign KJI = ~kji;  //complement 
assign KJJ = ~kjj;  //complement 
assign KJK = ~kjk;  //complement 
assign KJL = ~kjl;  //complement 
assign flm = ~FLM;  //complement 
assign fln = ~FLN;  //complement 
assign flo = ~FLO;  //complement 
assign flp = ~FLP;  //complement 
assign rbm = ~RBM;  //complement 
assign rbn = ~RBN;  //complement 
assign rbo = ~RBO;  //complement 
assign rbp = ~RBP;  //complement 
assign rcm = ~RCM;  //complement 
assign rcn = ~RCN;  //complement 
assign rco = ~RCO;  //complement 
assign rcp = ~RCP;  //complement 
assign ogi = ~OGI;  //complement 
assign ogj = ~OGJ;  //complement 
assign ogk = ~OGK;  //complement 
assign ogl = ~OGL;  //complement 
assign dbj =  bbg & cbh & cai  |  bbh & cai  |  bai  ; 
assign DBJ = ~dbj;  //complement 
assign fbc = ~FBC;  //complement 
assign fbi = ~FBI;  //complement 
assign QGG = ~qgg;  //complement 
assign QGH = ~qgh;  //complement 
assign QGI = ~qgi;  //complement 
assign QGJ = ~qgj;  //complement 
assign fcb = ~FCB;  //complement 
assign fce = ~FCE;  //complement 
assign fbd = ~FBD;  //complement 
assign fbj = ~FBJ;  //complement 
assign jab =  gaq & FAB  |  GAQ & fah  |  QGG  ; 
assign JAB = ~jab;  //complement 
assign jbb =  gaq & FAB  |  GAQ & fah  |  QGG  ; 
assign JBB = ~jbb; //complement 
assign ojc = ~OJC;  //complement 
assign qhc = ~QHC;  //complement 
assign fbe = ~FBE;  //complement 
assign fbk = ~FBK;  //complement 
assign gaa = ~GAA;  //complement 
assign gae = ~GAE;  //complement 
assign gak = ~GAK;  //complement 
assign gac = ~GAC;  //complement 
assign gai = ~GAI;  //complement 
assign gam = ~GAM;  //complement 
assign fbf = ~FBF;  //complement 
assign fbl = ~FBL;  //complement 
assign gag = ~GAG;  //complement 
assign gal = ~GAL;  //complement 
assign gan = ~GAN;  //complement 
assign gah = ~GAH;  //complement 
assign gaj = ~GAJ;  //complement 
assign gao = ~GAO;  //complement 
assign fca = ~FCA;  //complement 
assign fcd = ~FCD;  //complement 
assign gab = ~GAB;  //complement 
assign gad = ~GAD;  //complement 
assign gaf = ~GAF;  //complement 
assign qjm = ~QJM;  //complement 
assign oha = ~OHA;  //complement 
assign ECG =  BAM & BAN & BAO  ; 
assign ecg = ~ECG;  //complement 
assign ECH =  BAM & BAN & BAO  ; 
assign ech = ~ECH;  //complement 
assign ogm = ~OGM;  //complement 
assign ogn = ~OGN;  //complement 
assign ogo = ~OGO;  //complement 
assign ogp = ~OGP;  //complement 
assign fcc = ~FCC;  //complement 
assign fcf = ~FCF;  //complement 
assign ECA =  BAM & cam  ; 
assign eca = ~ECA;  //complement 
assign ECB =  BAN & can  ; 
assign ecb = ~ECB;  //complement 
assign ECC =  BAO & cao  ; 
assign ecc = ~ECC;  //complement 
assign dbk =  bbg & cbh & cai & caj  |  bbh & cai & caj  |  bai & caj  |  baj  ; 
assign DBK = ~dbk;  //complement 
assign bbi = ~BBI;  //complement 
assign bai = ~BAI;  //complement 
assign CAI = ~cai;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign dbl =  bbg & cbh & cai & caj & cak  |  bbh & cai & caj & cak  |  bai & caj & cak  |  baj & cak  |  bak  ; 
assign DBL = ~dbl;  //complement 
assign DBD =  CBG & BBH & BAI  |  CBH & BAI  |  CAI  ; 
assign dbd = ~DBD;  //complement 
assign baj = ~BAJ;  //complement 
assign CAJ = ~caj;  //complement 
assign AHI = ~ahi;  //complement 
assign AHJ = ~ahj;  //complement 
assign AHK = ~ahk;  //complement 
assign AHL = ~ahl;  //complement 
assign EBC =  BBI & cai  ; 
assign ebc = ~EBC;  //complement 
assign EBD =  BAJ & caj  ; 
assign ebd = ~EBD;  //complement 
assign bao = ~BAO;  //complement 
assign CAO = ~cao;  //complement 
assign bak = ~BAK;  //complement 
assign CAK = ~cak;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign EBE =  BAK & cak  ; 
assign ebe = ~EBE;  //complement 
assign EBF =  BAL & cal  ; 
assign ebf = ~EBF;  //complement 
assign DBG =  CBG & BBH & BAI & BAJ & BAK & BAL  |  CBH & BAI & BAJ & BAK & BAL  |  CAI & BAJ & BAK & BAL  |  CAJ & BAK & BAL  |  CAK & BAL  |  CAL  ; 
assign dbg = ~DBG;  //complement 
assign bal = ~BAL;  //complement 
assign CAL = ~cal;  //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign EBG =  BAG & BAH & BAI & BAJ & BAK & BAL  ; 
assign ebg = ~EBG;  //complement  
assign jea =  qdf & qdg & qec & qed  ; 
assign JEA = ~jea;  //complement 
assign DBF =  CBG & BBH & BAI & BAJ & BAK  |  CBH & BAI & BAJ & BAK  |  CAI & BAJ & BAK  |  CAJ & BAK  |  CAK  ; 
assign dbf = ~DBF;  //complement 
assign bam = ~BAM;  //complement 
assign CAM = ~cam;  //complement 
assign AHM = ~ahm;  //complement 
assign AHN = ~ahn;  //complement 
assign AHO = ~aho;  //complement 
assign dce =  bam  ; 
assign DCE = ~dce;  //complement 
assign dcf =  can & bam  |  ban  ; 
assign DCF = ~dcf;  //complement 
assign DCD =  CAM & BAN & BAO  |  CAN & BAO  |  CAO  ; 
assign dcd = ~DCD;  //complement 
assign ban = ~BAN;  //complement 
assign CAN = ~can;  //complement 
assign ado = ~ADO;  //complement 
assign dcb = ~DCB;  //complement 
assign dcc = ~DCC;  //complement 
assign bbg = ~BBG;  //complement 
assign CBG = ~cbg;  //complement 
assign DBE =  CBG & BBH & BAI & BAJ  |  CBH & BAI & BAJ  |  CAI & BAJ  |  CAJ  ; 
assign dbe = ~DBE;  //complement 
assign adp = ~ADP;  //complement 
assign QJA = ~qja;  //complement 
assign bbh = ~BBH;  //complement 
assign CBH = ~cbh;  //complement 
assign tda = ~TDA;  //complement 
assign tdb = ~TDB;  //complement 
assign tdc = ~TDC;  //complement 
assign tdd = ~TDD;  //complement 
assign AHP = ~ahp;  //complement 
assign rba = ~RBA;  //complement 
assign rbb = ~RBB;  //complement 
assign rbc = ~RBC;  //complement 
assign rbd = ~RBD;  //complement 
assign rca = ~RCA;  //complement 
assign rcb = ~RCB;  //complement 
assign rcc = ~RCC;  //complement 
assign rcd = ~RCD;  //complement 
assign QFB = ~qfb;  //complement 
assign raa = ~RAA;  //complement 
assign rab = ~RAB;  //complement 
assign qec = ~QEC;  //complement 
assign qef = ~QEF;  //complement 
assign qeg = ~QEG;  //complement 
assign qeh = ~QEH;  //complement 
assign KJA = ~kja;  //complement 
assign KJB = ~kjb;  //complement 
assign KJC = ~kjc;  //complement 
assign KJD = ~kjd;  //complement 
assign rac = ~RAC;  //complement 
assign rad = ~RAD;  //complement 
assign fla = ~FLA;  //complement 
assign flb = ~FLB;  //complement 
assign flc = ~FLC;  //complement 
assign fld = ~FLD;  //complement 
assign KKA = ~kka;  //complement 
assign KKB = ~kkb;  //complement 
assign KKC = ~kkc;  //complement 
assign KKD = ~kkd;  //complement 
assign QFC = ~qfc;  //complement 
assign fpa = ~FPA;  //complement 
assign fpb = ~FPB;  //complement 
assign fpc = ~FPC;  //complement 
assign fpd = ~FPD;  //complement 
assign KKE = ~kke;  //complement 
assign KKF = ~kkf;  //complement 
assign KKG = ~kkg;  //complement 
assign KKH = ~kkh;  //complement 
assign qga = ~QGA;  //complement 
assign qgb = ~QGB;  //complement 
assign fpe = ~FPE;  //complement 
assign fpf = ~FPF;  //complement 
assign fpg = ~FPG;  //complement 
assign fph = ~FPH;  //complement 
assign KJE = ~kje;  //complement 
assign KJF = ~kjf;  //complement 
assign KJG = ~kjg;  //complement 
assign KJH = ~kjh;  //complement 
assign rae = ~RAE;  //complement 
assign raf = ~RAF;  //complement 
assign fle = ~FLE;  //complement 
assign flf = ~FLF;  //complement 
assign flg = ~FLG;  //complement 
assign flh = ~FLH;  //complement 
assign QFA = ~qfa;  //complement 
assign rag = ~RAG;  //complement 
assign rah = ~RAH;  //complement 
assign qea = ~QEA;  //complement 
assign qeb = ~QEB;  //complement 
assign qed = ~QED;  //complement 
assign qee = ~QEE;  //complement 
assign TBA = ~tba;  //complement 
assign rbe = ~RBE;  //complement 
assign rbf = ~RBF;  //complement 
assign rbg = ~RBG;  //complement 
assign rbh = ~RBH;  //complement 
assign rce = ~RCE;  //complement 
assign rcf = ~RCF;  //complement 
assign rcg = ~RCG;  //complement 
assign rch = ~RCH;  //complement 
assign oga = ~OGA;  //complement 
assign ogb = ~OGB;  //complement 
assign ogc = ~OGC;  //complement 
assign ogd = ~OGD;  //complement 
assign daj =  baa & cab & cac  |  bab & cac  |  bac  ; 
assign DAJ = ~daj;  //complement 
assign faa = ~FAA;  //complement 
assign fag = ~FAG;  //complement 
assign dak =  bba & cbb & cac & cad  |  bbb & cac & cad  |  bac & cad  |  bad  ; 
assign DAK = ~dak;  //complement 
assign THA = gap; 
assign tha = ~THA; //complement 
assign THB = gap; 
assign thb = ~THB;  //complement 
assign THC = gap; 
assign thc = ~THC;  //complement 
assign THD = gap; 
assign thd = ~THD;  //complement 
assign fba = ~FBA;  //complement 
assign fbg = ~FBG;  //complement 
assign fab = ~FAB;  //complement 
assign fah = ~FAH;  //complement 
assign jca =  gaq & FAA  |  GAQ & fag  |  QGG  ; 
assign JCA = ~jca;  //complement 
assign jaa =  gaq & FAA  |  GAQ & fag  |  QGG  ; 
assign JAA = ~jaa; //complement 
assign jba =  gaq & FAA  |  GAQ & fag  |  QGG  ; 
assign JBA = ~jba;  //complement 
assign qya = ~QYA;  //complement 
assign oia = ~OIA;  //complement 
assign GCA = ~gca;  //complement 
assign GAP = ~gap;  //complement 
assign fae = ~FAE;  //complement 
assign fak = ~FAK;  //complement 
assign fad = ~FAD;  //complement 
assign GBA = ~gba;  //complement 
assign GAQ = ~gaq;  //complement 
assign faf = ~FAF;  //complement 
assign fal = ~FAL;  //complement 
assign oja = ~OJA;  //complement 
assign ojb = ~OJB;  //complement 
assign qha = ~QHA;  //complement 
assign qhb = ~QHB;  //complement 
assign bbc = ~BBC;  //complement 
assign fac = ~FAC;  //complement 
assign fai = ~FAI;  //complement 
assign qei = ~QEI;  //complement 
assign qej = ~QEJ;  //complement 
assign qek = ~QEK;  //complement 
assign faj = ~FAJ;  //complement 
assign oge = ~OGE;  //complement 
assign ogf = ~OGF;  //complement 
assign ogg = ~OGG;  //complement 
assign ogh = ~OGH;  //complement 
assign fbb = ~FBB;  //complement 
assign fbh = ~FBH;  //complement 
assign dbh =  bag  ; 
assign DBH = ~dbh;  //complement 
assign dbi =  cah & bag  |  bah  ; 
assign DBI = ~dbi;  //complement 
assign dah =  baa  ; 
assign DAH = ~dah;  //complement 
assign dai =  cab & baa  |  bab  ; 
assign DAI = ~dai;  //complement 
assign bba = ~BBA;  //complement 
assign CBA = ~cba;  //complement 
assign baa = ~BAA;  //complement 
assign CAA = ~caa;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign dal =  bba & cbb & cac & cad & cae  |  bbb & cac & cad & cae  |  bac & cad & cae  |  bad & cae  |  bae  ; 
assign DAL = ~dal;  //complement 
assign bbb = ~BBB;  //complement 
assign CBB = ~cbb;  //complement 
assign bab = ~BAB;  //complement 
assign CAB = ~cab;  //complement 
assign AHA = ~aha;  //complement 
assign AHB = ~ahb;  //complement 
assign AHC = ~ahc;  //complement 
assign AHD = ~ahd;  //complement 
assign DAB =  CAA  ; 
assign dab = ~DAB;  //complement 
assign DAC =  BAB & CAA  |  CAB  ; 
assign dac = ~DAC;  //complement 
assign CAG = ~cag;  //complement 
assign bac = ~BAC;  //complement 
assign CAC = ~cac;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign EAG =  BAA & BAB & BBC & BAD & BAE & BAF  ; 
assign eag = ~EAG;  //complement  
assign DAG =  CBA & BBB & BAC & BAD & BAE & BAF  |  CBB & BAC & BAD & BAE & BAF  |  CAC & BAD & BAE & BAF  |  CAD & BAE & BAF  |  CAE & BAF  |  CAF  ; 
assign dag = ~DAG;  //complement 
assign bad = ~BAD;  //complement 
assign CAD = ~cad;  //complement 
assign ade = ~ADE;  //complement 
assign DAF =  CAA & BAB & BBC & BAD & BAE  |  CAB & BBC & BAD & BAE  |  CBC & BAD & BAE  |  CAD & BAE  |  CAE  ; 
assign daf = ~DAF;  //complement 
assign DDG =  CBA & BBB & BAC & BAD & BAE & BAF  |  CBB & BAC & BAD & BAE & BAF  |  CAC & BAD & BAE & BAF  |  CAD & BAE & BAF  |  CAE & BAF  |  CAF  ; 
assign ddg = ~DDG;  //complement 
assign bae = ~BAE;  //complement 
assign CAE = ~cae;  //complement 
assign adf = ~ADF;  //complement 
assign EAD =  BAD & cad  ; 
assign ead = ~EAD;  //complement 
assign EAE =  BAE & cae  ; 
assign eae = ~EAE;  //complement 
assign EAF =  BAF & caf  ; 
assign eaf = ~EAF;  //complement 
assign DAE =  CAA & BBB & BAC & BAD  |  CAB & BAC & BAD  |  CAC & BAD  |  CAD  ; 
assign dae = ~DAE;  //complement 
assign baf = ~BAF;  //complement 
assign CAF = ~caf;  //complement 
assign AHE = ~ahe;  //complement 
assign AHF = ~ahf;  //complement 
assign AHG = ~ahg;  //complement 
assign AHH = ~ahh;  //complement 
assign EAA =  BAA & caa  ; 
assign eaa = ~EAA;  //complement 
assign EAB =  BAB & cab  ; 
assign eab = ~EAB;  //complement 
assign EAC =  BBC & cbc  ; 
assign eac = ~EAC;  //complement 
assign DAD =  CAA & BBB & BAC  |  CAB & BAC  |  CAC  ; 
assign dad = ~DAD;  //complement 
assign bag = ~BAG;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign EBA =  BAG & cag  ; 
assign eba = ~EBA;  //complement 
assign EBB =  BAH & cah  ; 
assign ebb = ~EBB;  //complement 
assign DBB =  CAG  ; 
assign dbb = ~DBB;  //complement 
assign DBC =  BAH & CAG  |  CAH  ; 
assign dbc = ~DBC;  //complement 
assign bah = ~BAH;  //complement 
assign CAH = ~cah;  //complement 
assign tde = ~TDE;  //complement 
assign tdf = ~TDF;  //complement 
assign tdg = ~TDG;  //complement 
assign tdh = ~TDH;  //complement 
assign fki = ~FKI;  //complement 
assign fkk = ~FKK;  //complement 
assign fkl = ~FKL;  //complement 
assign fkj = ~FKJ;  //complement 
assign KFI = ~kfi;  //complement 
assign KFJ = ~kfj;  //complement 
assign KFK = ~kfk;  //complement 
assign KFL = ~kfl;  //complement 
assign foi = ~FOI;  //complement 
assign foj = ~FOJ;  //complement 
assign fok = ~FOK;  //complement 
assign fol = ~FOL;  //complement 
assign KFM = ~kfm;  //complement 
assign KFN = ~kfn;  //complement 
assign fom = ~FOM;  //complement 
assign fon = ~FON;  //complement 
assign foo = ~FOO;  //complement 
assign fop = ~FOP;  //complement 
assign KFO = ~kfo;  //complement 
assign KFP = ~kfp;  //complement 
assign fkm = ~FKM;  //complement 
assign fkn = ~FKN;  //complement 
assign fko = ~FKO;  //complement 
assign fkp = ~FKP;  //complement 
assign HCI =  FOI & gae  |  FKI & GAE  ; 
assign hci = ~HCI;  //complement 
assign HCJ =  FOJ & gae  |  FKJ & GAE  ; 
assign hcj = ~HCJ;  //complement 
assign kci = ~KCI;  //complement 
assign koi = ~KOI;  //complement 
assign kpi = ~KPI;  //complement 
assign OFI = ~ofi;  //complement 
assign OFJ = ~ofj;  //complement 
assign kcj = ~KCJ;  //complement 
assign koj = ~KOJ;  //complement 
assign kpj = ~KPJ;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign HCO =  FOO & gal  |  FKO & GAL  ; 
assign hco = ~HCO;  //complement 
assign HCP =  FOP & gal  |  FKP & GAL  ; 
assign hcp = ~HCP;  //complement 
assign HCK =  FOK & gak  |  FKK & GAK  ; 
assign hck = ~HCK;  //complement 
assign HCL =  FOL & gak  |  FKL & GAK  ; 
assign hcl = ~HCL;  //complement 
assign kck = ~KCK;  //complement 
assign kok = ~KOK;  //complement 
assign kpk = ~KPK;  //complement 
assign NCA = fca & ~GAP & ~GCA  |  fcd & ~GAP & GCA  |  FCA & GAP & ~GCA  |  FCD & GAP & GCA; 
assign nca = ~NCA;  //complement 
assign JDM =  tqa & QXL  |  tma & QXL  |  QXC  |  QXF  |  QXI  |  QXM  ;
assign jdm = ~JDM;  //complement 
assign OFK = ~ofk;  //complement 
assign OFL = ~ofl;  //complement 
assign kcl = ~KCL;  //complement 
assign kol = ~KOL;  //complement 
assign kpl = ~KPL;  //complement 
assign NBA = FBG & ~gan & ~gba  |  FBA & ~gan & gba  |  fbg & gan & ~gba  |  fba & gan & gba; 
assign nba = ~NBA;  //complement 
assign JDC =  QXA  |  QXD  |  QXG  |  QXJ  ; 
assign jdc = ~JDC;  //complement 
assign HCM =  FOM & gaj  |  FKM & GAJ  ; 
assign hcm = ~HCM;  //complement 
assign HCN =  FON & gaj  |  FKN & GAJ  ; 
assign hcn = ~HCN;  //complement 
assign kcm = ~KCM;  //complement 
assign kom = ~KOM;  //complement 
assign kpm = ~KPM;  //complement 
assign JDL =  QXC  |  QXF  |  QXI  |  QXL  ; 
assign jdl = ~JDL;  //complement 
assign OFM = ~ofm;  //complement 
assign OFN = ~ofn;  //complement 
assign kcn = ~KCN;  //complement 
assign kon = ~KON;  //complement 
assign CBC = ~cbc;  //complement 
assign kco = ~KCO;  //complement 
assign koo = ~KOO;  //complement 
assign JDA =  QXA  |  QXD  |  QXG  |  QXJ  ; 
assign jda = ~JDA;  //complement 
assign JDB =  QXA  |  QXD  |  QXG  |  QXJ  ; 
assign jdb = ~JDB; //complement 
assign OFO = ~ofo;  //complement 
assign OFP = ~ofp;  //complement 
assign kcp = ~KCP;  //complement 
assign kop = ~KOP;  //complement 
assign tof = ~TOF;  //complement 
assign tpf = ~TPF;  //complement 
assign LCI =  KOI & TQO  |  KCM & TRK  ; 
assign lci = ~LCI;  //complement 
assign LFI =  KOI & TQO  |  KCM & TRK  ; 
assign lfi = ~LFI; //complement 
assign LII =  KOI & TQO  |  KCM & TRK  ; 
assign lii = ~LII;  //complement 
assign OCI = ~oci;  //complement 
assign OKA = ~oka;  //complement 
assign QKJ = ~qkj;  //complement 
assign QKK = ~qkk;  //complement 
assign QKL = ~qkl;  //complement 
assign tmf = ~TMF;  //complement 
assign tnf = ~TNF;  //complement 
assign LCJ =  KOJ & TQK  |  KCN & TRK  ; 
assign lcj = ~LCJ;  //complement 
assign LFJ =  KOJ & TQK  |  KCN & TRK  ; 
assign lfj = ~LFJ; //complement 
assign OCJ = ~ocj;  //complement 
assign OCN = ~ocn;  //complement 
assign tqk = ~TQK;  //complement 
assign tql = ~TQL;  //complement 
assign trk = ~TRK;  //complement 
assign trl = ~TRL;  //complement 
assign LCK =  KOK & TQK  |  KCO & TRK  ; 
assign lck = ~LCK;  //complement 
assign LFK =  KOK & TQK  |  KCO & TRK  ; 
assign lfk = ~LFK; //complement 
assign OCK = ~ock;  //complement 
assign AGI = ~agi;  //complement 
assign AGJ = ~agj;  //complement 
assign AGK = ~agk;  //complement 
assign AGL = ~agl;  //complement 
assign tuj =  gam & FAE  |  GAM & fak  |  QGD  ; 
assign TUJ = ~tuj;  //complement 
assign tuk =  gam & FAE  |  GAM & fak  |  QGD  ; 
assign TUK = ~tuk; //complement 
assign tul =  gam & FAE  |  GAM & fak  |  QGD  ; 
assign TUL = ~tul;  //complement 
assign LCL =  KOL & TQK  |  KCP & TRK  ; 
assign lcl = ~LCL;  //complement 
assign LFL =  KOL & TQK  |  KCP & TRK  ; 
assign lfl = ~LFL; //complement 
assign OCL = ~ocl;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign tvj =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVJ = ~tvj;  //complement 
assign tvk =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVK = ~tvk; //complement 
assign tvl =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVL = ~tvl;  //complement 
assign LCM =  KOM & TQL  ; 
assign lcm = ~LCM;  //complement 
assign OCM = ~ocm;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign tsk = ~TSK;  //complement 
assign tsl = ~TSL;  //complement 
assign ttk = ~TTK;  //complement 
assign ttl = ~TTL;  //complement 
assign LCN =  KON & TQL  ; 
assign lcn = ~LCN;  //complement 
assign AGM = ~agm;  //complement 
assign AGN = ~agn;  //complement 
assign AGO = ~ago;  //complement 
assign AGP = ~agp;  //complement 
assign QKF = ~qkf;  //complement 
assign QKG = ~qkg;  //complement 
assign QKH = ~qkh;  //complement 
assign QKI = ~qki;  //complement 
assign LCO =  KOO & TQL  ; 
assign lco = ~LCO;  //complement 
assign OCO = ~oco;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign LCP =  KOP & TQL  ; 
assign lcp = ~LCP;  //complement 
assign LFP =  KOP & TQL  ; 
assign lfp = ~LFP; //complement 
assign OCP = ~ocp;  //complement 
assign tea = ~TEA;  //complement 
assign fka = ~FKA;  //complement 
assign fkb = ~FKB;  //complement 
assign fkc = ~FKC;  //complement 
assign fkd = ~FKD;  //complement 
assign KFB = ~kfb;  //complement 
assign KFC = ~kfc;  //complement 
assign KFD = ~kfd;  //complement 
assign foa = ~FOA;  //complement 
assign fob = ~FOB;  //complement 
assign foc = ~FOC;  //complement 
assign fod = ~FOD;  //complement 
assign KFE = ~kfe;  //complement 
assign KFF = ~kff;  //complement 
assign foe = ~FOE;  //complement 
assign fof = ~FOF;  //complement 
assign fog = ~FOG;  //complement 
assign foh = ~FOH;  //complement 
assign KFG = ~kfg;  //complement 
assign KFH = ~kfh;  //complement 
assign KFA = ~kfa;  //complement 
assign fke = ~FKE;  //complement 
assign fkf = ~FKF;  //complement 
assign fkg = ~FKG;  //complement 
assign fkh = ~FKH;  //complement 
assign HCA =  FOA & gae  |  FKA & GAE  ; 
assign hca = ~HCA;  //complement 
assign HCB =  FOB & gae  |  FKB & GAE  ; 
assign hcb = ~HCB;  //complement 
assign kca = ~KCA;  //complement 
assign koa = ~KOA;  //complement 
assign kpa = ~KPA;  //complement 
assign QBE = ~qbe;  //complement 
assign QBH = ~qbh;  //complement 
assign OFA = ~ofa;  //complement 
assign OFB = ~ofb;  //complement 
assign kcb = ~KCB;  //complement 
assign kob = ~KOB;  //complement 
assign kpb = ~KPB;  //complement 
assign QBF = ~qbf;  //complement 
assign QBG = ~qbg;  //complement 
assign HCC =  FOC & gak  |  FKC & GAK  ; 
assign hcc = ~HCC;  //complement 
assign HCD =  FOD & gak  |  FKD & GAK  ; 
assign hcd = ~HCD;  //complement 
assign kcc = ~KCC;  //complement 
assign koc = ~KOC;  //complement 
assign kpc = ~KPC;  //complement 
assign NCB = fcb & ~GAP & ~GCA  |  fce & ~GAP & GCA  |  FCB & GAP & ~GCA  |  FCE & GAP & GCA; 
assign ncb = ~NCB;  //complement 
assign qxj = ~QXJ;  //complement 
assign qxk = ~QXK;  //complement 
assign qxl = ~QXL;  //complement 
assign OFC = ~ofc;  //complement 
assign OFD = ~ofd;  //complement 
assign kcd = ~KCD;  //complement 
assign kod = ~KOD;  //complement 
assign kpd = ~KPD;  //complement 
assign NBB = FBH & ~gan & ~gba  |  FBB & ~gan & gba  |  fbh & gan & ~gba  |  fbb & gan & gba; 
assign nbb = ~NBB;  //complement 
assign QXA = ~qxa;  //complement 
assign QXB = ~qxb;  //complement 
assign QXC = ~qxc;  //complement 
assign HCE =  FOE & gaj  |  FKE & GAJ  ; 
assign hce = ~HCE;  //complement 
assign HCF =  FOF & gaj  |  FKF & GAJ  ; 
assign hcf = ~HCF;  //complement 
assign kce = ~KCE;  //complement 
assign koe = ~KOE;  //complement 
assign kpe = ~KPE;  //complement 
assign QBA = ~qba;  //complement 
assign QBB = ~qbb;  //complement 
assign LCC =  KOC & TQI  |  KCG & TRI  |  KOK & TSI  |  KCO & TTI  ; 
assign lcc = ~LCC;  //complement 
assign OFE = ~ofe;  //complement 
assign OFF = ~off;  //complement 
assign kcf = ~KCF;  //complement 
assign kof = ~KOF;  //complement 
assign QBC = ~qbc;  //complement 
assign QBD = ~qbd;  //complement 
assign HCG =  FOG & gal  |  FKG & GAL  ; 
assign hcg = ~HCG;  //complement 
assign HCH =  FOH & gal  |  FKH & GAL  ; 
assign hch = ~HCH;  //complement 
assign kcg = ~KCG;  //complement 
assign kog = ~KOG;  //complement 
assign OFG = ~ofg;  //complement 
assign OFH = ~ofh;  //complement 
assign kch = ~KCH;  //complement 
assign koh = ~KOH;  //complement 
assign toe = ~TOE;  //complement 
assign tpe = ~TPE;  //complement 
assign LCA =  KOA & TQM  |  KCE & TRI  |  KOI & TSK  |  KPM & TTI  ; 
assign lca = ~LCA;  //complement 
assign LFA =  KOA & TQM  |  KCE & TRI  |  KOI & TSK  |  KPM & TTI  ; 
assign lfa = ~LFA; //complement 
assign LIA =  KOA & TQM  |  KCE & TRI  |  KOI & TSK  |  KPM & TTI  ; 
assign lia = ~LIA;  //complement 
assign OCA = ~oca;  //complement 
assign QAC = ~qac;  //complement 
assign QAD = ~qad;  //complement 
assign QAE = ~qae;  //complement 
assign tme = ~TME;  //complement 
assign tne = ~TNE;  //complement 
assign LCB =  KOB & TQI  |  KCF & TRI  |  KOJ & TSI  |  KCN & TTI  ; 
assign lcb = ~LCB;  //complement 
assign LFB =  KOB & TQI  |  KCF & TRI  |  KOJ & TSI  |  KCN & TTI  ; 
assign lfb = ~LFB; //complement 
assign OCB = ~ocb;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign tqi = ~TQI;  //complement 
assign tqj = ~TQJ;  //complement 
assign tri = ~TRI;  //complement 
assign trj = ~TRJ;  //complement 
assign OCG = ~ocg;  //complement 
assign OCC = ~occ;  //complement 
assign AGA = ~aga;  //complement 
assign AGB = ~agb;  //complement 
assign AGC = ~agc;  //complement 
assign AGD = ~agd;  //complement 
assign jac =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JAC = ~jac;  //complement 
assign jbc =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JBC = ~jbc; //complement 
assign jcc =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JCC = ~jcc;  //complement 
assign LCD =  KOD & TQI  |  KCH & TRI  |  KOL & TSI  |  KCP & TTI  ; 
assign lcd = ~LCD;  //complement 
assign LFD =  KOD & TQI  |  KCH & TRI  |  KOL & TSI  |  KCP & TTI  ; 
assign lfd = ~LFD; //complement 
assign OCD = ~ocd;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign jfc =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JFC = ~jfc;  //complement 
assign jhc =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JHC = ~jhc; //complement 
assign LCE =  KOE & TQJ  |  KCI & TRJ  |  KOM & TSJ  ; 
assign lce = ~LCE;  //complement 
assign OCE = ~oce;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign tsi = ~TSI;  //complement 
assign tsj = ~TSJ;  //complement 
assign tti = ~TTI;  //complement 
assign ttj = ~TTJ;  //complement 
assign LCF =  KOF & TQJ  |  KCJ & TRJ  |  KON & TSJ  ; 
assign lcf = ~LCF;  //complement 
assign OCF = ~ocf;  //complement 
assign AGE = ~age;  //complement 
assign AGF = ~agf;  //complement 
assign AGG = ~agg;  //complement 
assign AGH = ~agh;  //complement 
assign jad =  gai & FAD  |  GAI & faj  |  QGF  ; 
assign JAD = ~jad;  //complement 
assign jbd =  gai & FAD  |  GAI & faj  |  QGF  ; 
assign JBD = ~jbd; //complement 
assign jcd =  gai & FAD  |  GAI & faj  |  QGF  ; 
assign JCD = ~jcd;  //complement 
assign LCG =  KOG & TQJ  |  KCK & TRJ  |  KOO & TSJ  ; 
assign lcg = ~LCG;  //complement 
assign jgc =  gai & FAC  |  GAI & fai  |  QGF  ; 
assign JGC = ~jgc;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign TGE = ~tge;  //complement 
assign TGF = ~tgf;  //complement 
assign LCH =  KOH & TQJ  |  KCL & TRJ  |  KOP & TSJ  ; 
assign lch = ~LCH;  //complement 
assign LFH =  KOH & TQJ  |  KCL & TRJ  |  KOP & TSJ  ; 
assign lfh = ~LFH; //complement 
assign OCH = ~och;  //complement 
assign QAA = ~qaa;  //complement 
assign QAB = ~qab;  //complement 
assign fji = ~FJI;  //complement 
assign fjj = ~FJJ;  //complement 
assign fjl = ~FJL;  //complement 
assign fjk = ~FJK;  //complement 
assign KEI = ~kei;  //complement 
assign KEK = ~kek;  //complement 
assign KEL = ~kel;  //complement 
assign fni = ~FNI;  //complement 
assign fnj = ~FNJ;  //complement 
assign fnk = ~FNK;  //complement 
assign fnl = ~FNL;  //complement 
assign fjn = ~FJN;  //complement 
assign fjp = ~FJP;  //complement 
assign KEM = ~kem;  //complement 
assign KEN = ~ken;  //complement 
assign fnm = ~FNM;  //complement 
assign fnn = ~FNN;  //complement 
assign fno = ~FNO;  //complement 
assign fnp = ~FNP;  //complement 
assign KEO = ~keo;  //complement 
assign KEP = ~kep;  //complement 
assign KEJ = ~kej;  //complement 
assign LFC =  KOC & TQI  |  KCG & TRI  |  KOK & TSI  |  KCO & TTI  ; 
assign lfc = ~LFC;  //complement 
assign fjm = ~FJM;  //complement 
assign fjo = ~FJO;  //complement 
assign HBI =  FNI & gae  |  FJI & GAE  ; 
assign hbi = ~HBI;  //complement 
assign HBJ =  FNJ & gae  |  FJJ & GAE  ; 
assign hbj = ~HBJ;  //complement 
assign kbi = ~KBI;  //complement 
assign kmi = ~KMI;  //complement 
assign kni = ~KNI;  //complement 
assign OEI = ~oei;  //complement 
assign OEJ = ~oej;  //complement 
assign kbj = ~KBJ;  //complement 
assign kmj = ~KMJ;  //complement 
assign knj = ~KNJ;  //complement 
assign HBL =  FNL & gag  |  FJL & GAG  ; 
assign hbl = ~HBL;  //complement 
assign kbk = ~KBK;  //complement 
assign kmk = ~KMK;  //complement 
assign knk = ~KNK;  //complement 
assign NCC = fcc & ~GAP & ~GCA  |  fcf & ~GAP & GCA  |  FCC & GAP & ~GCA  |  FCF & GAP & GCA; 
assign ncc = ~NCC;  //complement 
assign QXD = ~qxd;  //complement 
assign QXE = ~qxe;  //complement 
assign QXF = ~qxf;  //complement 
assign OEK = ~oek;  //complement 
assign OEL = ~oel;  //complement 
assign kbl = ~KBL;  //complement 
assign kml = ~KML;  //complement 
assign knl = ~KNL;  //complement 
assign NBC = FBI & ~gan & ~gba  |  FBC & ~gan & gba  |  fbi & gan & ~gba  |  fbc & gan & gba; 
assign nbc = ~NBC;  //complement 
assign JDD =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jdd = ~JDD;  //complement 
assign JDE =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jde = ~JDE; //complement 
assign JDF =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jdf = ~JDF;  //complement 
assign HBM =  FNM & gah  |  FJM & GAH  ; 
assign hbm = ~HBM;  //complement 
assign HBN =  FNN & gah  |  FJN & GAH  ; 
assign hbn = ~HBN;  //complement 
assign kbm = ~KBM;  //complement 
assign kmm = ~KMM;  //complement 
assign knm = ~KNM;  //complement 
assign OEM = ~oem;  //complement 
assign OEN = ~oen;  //complement 
assign kbn = ~KBN;  //complement 
assign kmn = ~KMN;  //complement 
assign HBO =  FNO & gaf  |  FJO & GAF  ; 
assign hbo = ~HBO;  //complement 
assign HBP =  FNP & gaf  |  FJP & GAF  ; 
assign hbp = ~HBP;  //complement 
assign kbo = ~KBO;  //complement 
assign kmo = ~KMO;  //complement 
assign hbk = ~HBK;  //complement 
assign OEO = ~oeo;  //complement 
assign OEP = ~oep;  //complement 
assign kbp = ~KBP;  //complement 
assign kmp = ~KMP;  //complement 
assign tod = ~TOD;  //complement 
assign tpd = ~TPD;  //complement 
assign LBI =  KMI & TQM  |  KBM & TRG  |  KOA & TSK  |  KPE & TTG  ; 
assign lbi = ~LBI;  //complement 
assign LEI =  KMI & TQM  |  KBM & TRG  |  KOA & TSK  |  KPE & TTG  ; 
assign lei = ~LEI; //complement 
assign LHT =  KMI & TQM  |  KBM & TRG  |  KOA & TSK  |  KPE & TTG  ; 
assign lht = ~LHT;  //complement 
assign OBI = ~obi;  //complement 
assign tmd = ~TMD;  //complement 
assign tnd = ~TND;  //complement 
assign LBJ =  KMJ & TQG  |  KBN & TRG  |  KOB & TSG  |  KCF & TTG  ; 
assign lbj = ~LBJ;  //complement 
assign LEJ =  KMJ & TQG  |  KBN & TRG  |  KOB & TSG  |  KCF & TTG  ; 
assign lej = ~LEJ; //complement 
assign OBJ = ~obj;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign tqg = ~TQG;  //complement 
assign tqh = ~TQH;  //complement 
assign trg = ~TRG;  //complement 
assign trh = ~TRH;  //complement 
assign LBK =  KMK & TQG  |  KBO & TRG  |  KOC & TSG  |  KCG & TTG  ; 
assign lbk = ~LBK;  //complement 
assign LEK =  KMK & TQG  |  KBO & TRG  |  KOC & TSG  |  KCG & TTG  ; 
assign lek = ~LEK; //complement 
assign OBK = ~obk;  //complement 
assign AFI = ~afi;  //complement 
assign AFJ = ~afj;  //complement 
assign AFK = ~afk;  //complement 
assign AFL = ~afl;  //complement 
assign tug =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUG = ~tug;  //complement 
assign tuh =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUH = ~tuh; //complement 
assign tui =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUI = ~tui;  //complement 
assign LBL =  KML & TQG  |  KBP & TRG  |  KOD & TSG  |  KCH & TTG  ; 
assign lbl = ~LBL;  //complement 
assign LEL =  KML & TQG  |  KBP & TRG  |  KOD & TSG  |  KCH & TTG  ; 
assign lel = ~LEL; //complement 
assign OBL = ~obl;  //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign tvg =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVG = ~tvg;  //complement 
assign tvh =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVH = ~tvh; //complement 
assign tvi =  gao & FAF  |  QGE  |  GAO & fal  ; 
assign TVI = ~tvi;  //complement 
assign LBM =  KMM & TQH  |  KCA & TRH  |  KOE & TSH  |  KPI & TTH  ; 
assign lbm = ~LBM;  //complement 
assign OBM = ~obm;  //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign tsg = ~TSG;  //complement 
assign tsh = ~TSH;  //complement 
assign ttg = ~TTG;  //complement 
assign tth = ~TTH;  //complement 
assign LBN =  KMN & TQH  |  KCB & TRH  |  KOF & TSH  |  KPJ & TTH  ; 
assign lbn = ~LBN;  //complement 
assign OBN = ~obn;  //complement 
assign AFM = ~afm;  //complement 
assign AFN = ~afn;  //complement 
assign AFO = ~afo;  //complement 
assign AFP = ~afp;  //complement 
assign QKA = ~qka;  //complement 
assign QKD = ~qkd;  //complement 
assign QKE = ~qke;  //complement 
assign LBO =  KMO & TQH  |  KCC & TRH  |  KOG & TSH  |  KPK & TTH  ; 
assign lbo = ~LBO;  //complement 
assign OBO = ~obo;  //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign QKB = ~qkb;  //complement 
assign qkc = ~QKC;  //complement 
assign LBP =  KMP & TQH  |  KCD & TRH  |  KOH & TSH  |  KPL & TTH  ; 
assign lbp = ~LBP;  //complement 
assign LEP =  KMP & TQH  |  KCD & TRH  |  KOH & TSH  |  KPL & TTH  ; 
assign lep = ~LEP; //complement 
assign OBP = ~obp;  //complement 
assign qia = ~QIA;  //complement 
assign qib = ~QIB;  //complement 
assign fja = ~FJA;  //complement 
assign fjb = ~FJB;  //complement 
assign fjc = ~FJC;  //complement 
assign fjd = ~FJD;  //complement 
assign KEA = ~kea;  //complement 
assign KEB = ~keb;  //complement 
assign KEC = ~kec;  //complement 
assign KED = ~ked;  //complement 
assign fna = ~FNA;  //complement 
assign fnb = ~FNB;  //complement 
assign fnc = ~FNC;  //complement 
assign fnd = ~FND;  //complement 
assign KEE = ~kee;  //complement 
assign KEF = ~kef;  //complement 
assign fne = ~FNE;  //complement 
assign fnf = ~FNF;  //complement 
assign fng = ~FNG;  //complement 
assign fnh = ~FNH;  //complement 
assign KEG = ~keg;  //complement 
assign KEH = ~keh;  //complement 
assign fje = ~FJE;  //complement 
assign fjf = ~FJF;  //complement 
assign fjg = ~FJG;  //complement 
assign fjh = ~FJH;  //complement 
assign HBA =  FNA & gae  |  FJA & GAE  ; 
assign hba = ~HBA;  //complement 
assign HBB =  FNB & gae  |  FJB & GAE  ; 
assign hbb = ~HBB;  //complement 
assign kba = ~KBA;  //complement 
assign kma = ~KMA;  //complement 
assign kna = ~KNA;  //complement 
assign OEA = ~oea;  //complement 
assign OEB = ~oeb;  //complement 
assign kbb = ~KBB;  //complement 
assign kmb = ~KMB;  //complement 
assign knb = ~KNB;  //complement 
assign OEE = ~oee;  //complement 
assign HBC =  FNC & gag  |  FJC & GAG  ; 
assign hbc = ~HBC;  //complement 
assign HBD =  FND & gag  |  FJD & GAG  ; 
assign hbd = ~HBD;  //complement 
assign kbc = ~KBC;  //complement 
assign kmc = ~KMC;  //complement 
assign knc = ~KNC;  //complement 
assign QXM = ~qxm;  //complement 
assign OEC = ~oec;  //complement 
assign OED = ~oed;  //complement 
assign kbd = ~KBD;  //complement 
assign kmd = ~KMD;  //complement 
assign knd = ~KND;  //complement 
assign NBD = FBJ & ~gan & ~gba  |  FBD & ~gan & gba  |  fbj & gan & ~gba  |  fbd & gan & gba; 
assign nbd = ~NBD;  //complement 
assign JDG =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jdg = ~JDG;  //complement 
assign JDH =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jdh = ~JDH; //complement 
assign JDI =  QXB  |  QXE  |  QXK  |  QXH  ; 
assign jdi = ~JDI;  //complement 
assign HBE =  FNE & gah  |  FJE & GAH  ; 
assign hbe = ~HBE;  //complement 
assign HBF =  FNF & gah  |  FJF & GAH  ; 
assign hbf = ~HBF;  //complement 
assign kbe = ~KBE;  //complement 
assign kme = ~KME;  //complement 
assign kne = ~KNE;  //complement 
assign OEF = ~oef;  //complement 
assign kbf = ~KBF;  //complement 
assign kmf = ~KMF;  //complement 
assign HBG =  FNG & gaf  |  FJG & GAF  ; 
assign hbg = ~HBG;  //complement 
assign HBH =  FNH & gaf  |  FJH & GAF  ; 
assign hbh = ~HBH;  //complement 
assign kbg = ~KBG;  //complement 
assign kmg = ~KMG;  //complement 
assign OEG = ~oeg;  //complement 
assign OEH = ~oeh;  //complement 
assign kbh = ~KBH;  //complement 
assign kmh = ~KMH;  //complement 
assign toc = ~TOC;  //complement 
assign tpc = ~TPC;  //complement 
assign LBA =  KMA & TQN  |  KBE & TRE  |  KMI & TSL  |  KNM & TTE  ; 
assign lba = ~LBA;  //complement 
assign LEA =  KMA & TQN  |  KBE & TRE  |  KMI & TSL  |  KNM & TTE  ; 
assign lea = ~LEA; //complement 
assign LHA =  KMA & TQN  |  KBE & TRE  |  KMI & TSL  |  KNM & TTE  ; 
assign lha = ~LHA;  //complement 
assign OBA = ~oba;  //complement 
assign LAR =  KAQ & TQE  |  KAR & TQE  |  KLD & TRL  |  KLH & TSE  |  KQL & TTL  ;
assign lar = ~LAR;  //complement 
assign tmc = ~TMC;  //complement 
assign tnc = ~TNC;  //complement 
assign LBB =  KMB & TQE  |  KBF & TRE  |  KMJ & TSE  |  KBN & TTE  ; 
assign lbb = ~LBB;  //complement 
assign LEB =  KMB & TQE  |  KBF & TRE  |  KMJ & TSE  |  KBN & TTE  ; 
assign leb = ~LEB; //complement 
assign OBB = ~obb;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign tqe = ~TQE;  //complement 
assign tqf = ~TQF;  //complement 
assign tre = ~TRE;  //complement 
assign trf = ~TRF;  //complement 
assign LBC =  KMC & TQE  |  KBG & TRE  |  KMK & TSE  |  KBO & TTE  ; 
assign lbc = ~LBC;  //complement 
assign LEC =  KMC & TQE  |  KBG & TRE  |  KMK & TSE  |  KBO & TTE  ; 
assign lec = ~LEC; //complement 
assign OBC = ~obc;  //complement 
assign AFA = ~afa;  //complement 
assign AFB = ~afb;  //complement 
assign AFC = ~afc;  //complement 
assign AFD = ~afd;  //complement 
assign tud =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUD = ~tud;  //complement 
assign tue =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUE = ~tue; //complement 
assign tuf =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUF = ~tuf;  //complement 
assign LBD =  KMD & TQE  |  KBH & TRE  |  KML & TSE  |  KBP & TTE  ; 
assign lbd = ~LBD;  //complement 
assign LED =  KMD & TQE  |  KBH & TRE  |  KML & TSE  |  KBP & TTE  ; 
assign led = ~LED; //complement 
assign OBD = ~obd;  //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign tvd =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVD = ~tvd;  //complement 
assign tve =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVE = ~tve; //complement 
assign tvf =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVF = ~tvf;  //complement 
assign LBE =  KME & TQF  |  KBI & TRF  |  KMM & TSF  |  KPA & TTF  ; 
assign lbe = ~LBE;  //complement 
assign OBE = ~obe;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign tse = ~TSE;  //complement 
assign tsf = ~TSF;  //complement 
assign tte = ~TTE;  //complement 
assign ttf = ~TTF;  //complement 
assign LBF =  KMF & TQF  |  KBJ & TRF  |  KMN & TSF  |  KPB & TTF  ; 
assign lbf = ~LBF;  //complement 
assign OBF = ~obf;  //complement 
assign AFE = ~afe;  //complement 
assign AFF = ~aff;  //complement 
assign AFG = ~afg;  //complement 
assign AFH = ~afh;  //complement 
assign LBG =  KMG & TQF  |  KBK & TRF  |  KMO & TSF  |  KPC & TTF  ; 
assign lbg = ~LBG;  //complement 
assign OBG = ~obg;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign TGC = ~tgc;  //complement 
assign TGD = ~tgd;  //complement 
assign LBH =  KMH & TQF  |  KBL & TRF  |  KMP & TSF  |  KPD & TTF  ; 
assign lbh = ~LBH;  //complement 
assign LEH =  KMH & TQF  |  KBL & TRF  |  KMP & TSF  |  KPD & TTF  ; 
assign leh = ~LEH; //complement 
assign OBH = ~obh;  //complement 
assign fii = ~FII;  //complement 
assign fij = ~FIJ;  //complement 
assign fik = ~FIK;  //complement 
assign fil = ~FIL;  //complement 
assign KDI = ~kdi;  //complement 
assign KDJ = ~kdj;  //complement 
assign KDK = ~kdk;  //complement 
assign KDL = ~kdl;  //complement 
assign fmi = ~FMI;  //complement 
assign fmj = ~FMJ;  //complement 
assign fmk = ~FMK;  //complement 
assign fml = ~FML;  //complement 
assign KDM = ~kdm;  //complement 
assign KDN = ~kdn;  //complement 
assign fmm = ~FMM;  //complement 
assign fmn = ~FMN;  //complement 
assign fmo = ~FMO;  //complement 
assign fmp = ~FMP;  //complement 
assign KDO = ~kdo;  //complement 
assign KDP = ~kdp;  //complement 
assign fim = ~FIM;  //complement 
assign fin = ~FIN;  //complement 
assign fio = ~FIO;  //complement 
assign fip = ~FIP;  //complement 
assign HAI =  FMI & gaa  |  FII & GAA  ; 
assign hai = ~HAI;  //complement 
assign HAJ =  FMJ & gaa  |  FIJ & GAA  ; 
assign haj = ~HAJ;  //complement 
assign kai = ~KAI;  //complement 
assign kli = ~KLI;  //complement 
assign ODI = ~odi;  //complement 
assign ODJ = ~odj;  //complement 
assign kaj = ~KAJ;  //complement 
assign klj = ~KLJ;  //complement 
assign ODO = ~odo;  //complement 
assign HAK =  FMK & gac  |  FIK & GAC  ; 
assign hak = ~HAK;  //complement 
assign HAL =  FML & gac  |  FIL & GAC  ; 
assign hal = ~HAL;  //complement 
assign kak = ~KAK;  //complement 
assign klk = ~KLK;  //complement 
assign ODN = ~odn;  //complement 
assign NBF = fbf & ~GAN & ~GBA  |  fbl & ~GAN & GBA  |  FBF & GAN & ~GBA  |  FBL & GAN & GBA; 
assign nbf = ~NBF;  //complement 
assign ODK = ~odk;  //complement 
assign ODL = ~odl;  //complement 
assign kal = ~KAL;  //complement 
assign kll = ~KLL;  //complement 
assign kql = ~KQL;  //complement 
assign NBE = fbe & ~GAN & ~GBA  |  fbk & ~GAN & GBA  |  FBE & GAN & ~GBA  |  FBK & GAN & GBA; 
assign nbe = ~NBE;  //complement 
assign QXG = ~qxg;  //complement 
assign QXH = ~qxh;  //complement 
assign QXI = ~qxi;  //complement 
assign HAM =  FMM & gab  |  FIM & GAB  ; 
assign ham = ~HAM;  //complement 
assign HAN =  FMN & gab  |  FIN & GAB  ; 
assign han = ~HAN;  //complement 
assign kam = ~KAM;  //complement 
assign klm = ~KLM;  //complement 
assign kqm = ~KQM;  //complement 
assign ODM = ~odm;  //complement 
assign kln = ~KLN;  //complement 
assign HAO =  FMO & gad  |  FIO & GAD  ; 
assign hao = ~HAO;  //complement 
assign HAP =  FMP & gad  |  FIP & GAD  ; 
assign hap = ~HAP;  //complement 
assign kao = ~KAO;  //complement 
assign klo = ~KLO;  //complement 
assign kan = ~KAN;  //complement 
assign ODP = ~odp;  //complement 
assign kap = ~KAP;  //complement 
assign klp = ~KLP;  //complement 
assign tob = ~TOB;  //complement 
assign tpb = ~TPB;  //complement 
assign LAI =  KLI & TQN  |  KAM & TRC  |  KMA & TSL  |  KNE & TTC  ; 
assign lai = ~LAI;  //complement 
assign LDI =  KLI & TQN  |  KAM & TRC  |  KMA & TSL  |  KNE & TTC  ; 
assign ldi = ~LDI; //complement 
assign LGI =  KLI & TQN  |  KAM & TRC  |  KMA & TSL  |  KNE & TTC  ; 
assign lgi = ~LGI;  //complement 
assign OAI = ~oai;  //complement 
assign OAR = ~oar;  //complement 
assign tmb = ~TMB;  //complement 
assign tnb = ~TNB;  //complement 
assign LAJ =  KLJ & TQC  |  KAN & TRC  |  KMB & TSC  |  KBF & TTC  ; 
assign laj = ~LAJ;  //complement 
assign LDJ =  KLJ & TQC  |  KAN & TRC  |  KMB & TSC  |  KBF & TTC  ; 
assign ldj = ~LDJ; //complement 
assign OAJ = ~oaj;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign tqc = ~TQC;  //complement 
assign tqd = ~TQD;  //complement 
assign trc = ~TRC;  //complement 
assign trd = ~TRD;  //complement 
assign OAO = ~oao;  //complement 
assign OAK = ~oak;  //complement 
assign AEI = ~aei;  //complement 
assign AEJ = ~aej;  //complement 
assign AEK = ~aek;  //complement 
assign AEL = ~ael;  //complement 
assign qgc = ~QGC;  //complement 
assign qgd = ~QGD;  //complement 
assign qge = ~QGE;  //complement 
assign qgf = ~QGF;  //complement 
assign LAL =  KLL & TQC  |  KAP & TRC  |  KMD & TSC  |  KBH & TTC  ; 
assign lal = ~LAL;  //complement 
assign LDL =  KLL & TQC  |  KAP & TRC  |  KMD & TSC  |  KBH & TTC  ; 
assign ldl = ~LDL; //complement 
assign OAL = ~oal;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign TQM = ~tqm;  //complement 
assign TQN = ~tqn;  //complement 
assign TQO = ~tqo;  //complement 
assign LAM =  KLM & TQD  |  KBA & TRD  |  KME & TSD  |  KNI & TTD  ; 
assign lam = ~LAM;  //complement 
assign OAM = ~oam;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign tsc = ~TSC;  //complement 
assign tsd = ~TSD;  //complement 
assign ttc = ~TTC;  //complement 
assign ttd = ~TTD;  //complement 
assign LAN =  KLN & TQD  |  KBB & TRD  |  KMF & TSD  |  KNJ & TTD  ; 
assign lan = ~LAN;  //complement 
assign OAN = ~oan;  //complement 
assign AEM = ~aem;  //complement 
assign AEN = ~aen;  //complement 
assign AEO = ~aeo;  //complement 
assign AEP = ~aep;  //complement 
assign KAR = ~kar;  //complement 
assign LAO =  KLO & TQD  |  KBC & TRD  |  KMG & TSD  |  KNK & TTD  ; 
assign lao = ~LAO;  //complement 
assign LDO =  KLO & TQD  |  KBC & TRD  |  KMG & TSD  |  KNK & TTD  ; 
assign ldo = ~LDO; //complement 
assign LAK =  KLK & TQC  |  KAO & TRC  |  KMC & TSC  |  KBG & TTC  ; 
assign lak = ~LAK;  //complement 
assign LDK =  KLK & TQC  |  KAO & TRC  |  KMC & TSC  |  KBG & TTC  ; 
assign ldk = ~LDK; //complement 
assign aap = ~AAP;  //complement 
assign aao = ~AAO;  //complement 
assign kaq = ~KAQ;  //complement 
assign LAP =  KLP & TQD  |  KBD & TRD  |  KMH & TSD  |  KNL & TTD  ; 
assign lap = ~LAP;  //complement 
assign LDP =  KLP & TQD  |  KBD & TRD  |  KMH & TSD  |  KNL & TTD  ; 
assign ldp = ~LDP; //complement 
assign OAP = ~oap;  //complement 
assign QDI = ~qdi;  //complement 
assign kaa = ~KAA;  //complement 
assign qdc = ~QDC;  //complement 
assign qdf = ~QDF;  //complement 
assign qdg = ~QDG;  //complement 
assign kab = ~KAB;  //complement 
assign qdd = ~QDD;  //complement 
assign KDA = ~kda;  //complement 
assign KDB = ~kdb;  //complement 
assign fia = ~FIA;  //complement 
assign fib = ~FIB;  //complement 
assign fic = ~FIC;  //complement 
assign fid = ~FID;  //complement 
assign kac = ~KAC;  //complement 
assign kae = ~KAE;  //complement 
assign KDC = ~kdc;  //complement 
assign KDD = ~kdd;  //complement 
assign fma = ~FMA;  //complement 
assign fmb = ~FMB;  //complement 
assign fmc = ~FMC;  //complement 
assign fmd = ~FMD;  //complement 
assign kad = ~KAD;  //complement 
assign KDE = ~kde;  //complement 
assign KDF = ~kdf;  //complement 
assign fme = ~FME;  //complement 
assign fmf = ~FMF;  //complement 
assign fmg = ~FMG;  //complement 
assign fmh = ~FMH;  //complement 
assign KDG = ~kdg;  //complement 
assign KDH = ~kdh;  //complement 
assign fie = ~FIE;  //complement 
assign fif = ~FIF;  //complement 
assign fig = ~FIG;  //complement 
assign fih = ~FIH;  //complement 
assign qdh = ~QDH;  //complement 
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign qca = ~QCA;  //complement 
assign qcb = ~QCB;  //complement 
assign qcd = ~QCD;  //complement 
assign qce = ~QCE;  //complement 
assign qde = ~QDE;  //complement 
assign qci = ~QCI;  //complement 
assign qcc = ~QCC;  //complement 
assign qcf = ~QCF;  //complement 
assign qcg = ~QCG;  //complement 
assign qch = ~QCH;  //complement 
assign HAA =  FMA & gaa  |  FIA & GAA  ; 
assign haa = ~HAA;  //complement 
assign HAB =  FMB & gaa  |  FIB & GAA  ; 
assign hab = ~HAB;  //complement 
assign ODA = ~oda;  //complement 
assign ODB = ~odb;  //complement 
assign THE = gap; 
assign the = ~THE; //complement 
assign THF = gap; 
assign thf = ~THF;  //complement 
assign THG = gap; 
assign thg = ~THG;  //complement 
assign THH = gap; 
assign thh = ~THH;  //complement 
assign HAG =  FMG & gad  |  FIG & GAD  ; 
assign hag = ~HAG;  //complement 
assign HAH =  FMH & gad  |  FIH & GAD  ; 
assign hah = ~HAH;  //complement 
assign HAC =  FMC & gac  |  FIC & GAC  ; 
assign hac = ~HAC;  //complement 
assign HAD =  FMD & gac  |  FID & GAC  ; 
assign had = ~HAD;  //complement 
assign ODC = ~odc;  //complement 
assign ODD = ~odd;  //complement 
assign kld = ~KLD;  //complement 
assign JDJ =  QXC  |  QXF  |  QXI  |  QXL  ; 
assign jdj = ~JDJ;  //complement 
assign JDK =  QXC  |  QXF  |  QXI  |  QXL  ; 
assign jdk = ~JDK; //complement 
assign HAE =  FME & gab  |  FIE & GAB  ; 
assign hae = ~HAE;  //complement 
assign HAF =  FMF & gab  |  FIF & GAB  ; 
assign haf = ~HAF;  //complement 
assign ODE = ~ode;  //complement 
assign ODF = ~odf;  //complement 
assign kaf = ~KAF;  //complement 
assign QDJ = ~qdj;  //complement 
assign kag = ~KAG;  //complement 
assign jia =  qdb & qdj  ; 
assign JIA = ~jia;  //complement 
assign ODG = ~odg;  //complement 
assign ODH = ~odh;  //complement 
assign kah = ~KAH;  //complement 
assign klh = ~KLH;  //complement 
assign toa = ~TOA;  //complement 
assign tpa = ~TPA;  //complement 
assign LAA =  KAA & TQA  |  KAE & TRA  |  KLI & TSA  |  KQM & TTA  ; 
assign laa = ~LAA;  //complement 
assign OAA = ~oaa;  //complement 
assign TAA = ~taa;  //complement 
assign TAB = ~tab;  //complement 
assign TAC = ~tac;  //complement 
assign TAD = ~tad;  //complement 
assign tma = ~TMA;  //complement 
assign tna = ~TNA;  //complement 
assign LAB =  KAB & TQA  |  KAF & TRA  |  KLJ & TSA  |  KAN & TTA  ; 
assign lab = ~LAB;  //complement 
assign OAB = ~oab;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign tqa = ~TQA;  //complement 
assign tqb = ~TQB;  //complement 
assign tra = ~TRA;  //complement 
assign trb = ~TRB;  //complement 
assign OAG = ~oag;  //complement 
assign OAC = ~oac;  //complement 
assign AEA = ~aea;  //complement 
assign AEB = ~aeb;  //complement 
assign AEC = ~aec;  //complement 
assign AED = ~aed;  //complement 
assign tua =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUA = ~tua;  //complement 
assign tub =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUB = ~tub; //complement 
assign tuc =  gam & FAE  |  GAM & fak  |  QGC  ; 
assign TUC = ~tuc;  //complement 
assign LAD =  KAD & TQA  |  KAH & TRA  |  KLL & TSA  |  KAP & TTA  ; 
assign lad = ~LAD;  //complement 
assign LDD =  KAD & TQA  |  KAH & TRA  |  KLL & TSA  |  KAP & TTA  ; 
assign ldd = ~LDD; //complement 
assign OAD = ~oad;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign tva =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVA = ~tva;  //complement 
assign tvb =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVB = ~tvb; //complement 
assign tvc =  gao & FAF  |  QGD  |  GAO & fal  ; 
assign TVC = ~tvc;  //complement 
assign LAE =  KAE & TQB  |  KAI & TRB  |  KLM & TSB  |  KNA & TTB  ; 
assign lae = ~LAE;  //complement 
assign OAE = ~oae;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign tsa = ~TSA;  //complement 
assign tsb = ~TSB;  //complement 
assign tta = ~TTA;  //complement 
assign ttb = ~TTB;  //complement 
assign LAF =  KAF & TQB  |  KAJ & TRB  |  KLN & TSB  |  KNB & TTB  ; 
assign laf = ~LAF;  //complement 
assign OAF = ~oaf;  //complement 
assign AEE = ~aee;  //complement 
assign AEF = ~aef;  //complement 
assign AEG = ~aeg;  //complement 
assign AEH = ~aeh;  //complement 
assign LAG =  KAG & TQB  |  KAK & TRB  |  KLO & TSB  |  KNC & TTB  ; 
assign lag = ~LAG;  //complement 
assign LAC =  KAC & TQA  |  KAG & TRA  |  KLK & TSA  |  KAO & TTA  ; 
assign lac = ~LAC;  //complement 
assign LDC =  KAC & TQA  |  KAG & TRA  |  KLK & TSA  |  KAO & TTA  ; 
assign ldc = ~LDC; //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign TGA = ~tga;  //complement 
assign TGB = ~tgb;  //complement 
assign LAH =  KAH & TQB  |  KAL & TRB  |  KLP & TSB  |  KND & TTB  ; 
assign lah = ~LAH;  //complement 
assign LDH =  KAH & TQB  |  KAL & TRB  |  KLP & TSB  |  KND & TTB  ; 
assign ldh = ~LDH; //complement 
assign OAH = ~oah;  //complement 
assign TCA = ~tca;  //complement 
assign TCB = ~tcb;  //complement 
assign TCC = ~tcc;  //complement 
assign TCD = ~tcd;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iff = ~IFF; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
assign ihm = ~IHM; //complement 
assign ihn = ~IHN; //complement 
assign iho = ~IHO; //complement 
assign ihp = ~IHP; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ika = ~IKA; //complement 
assign ila = ~ILA; //complement 
always@(posedge IZZ )
   begin 
 RBI <= RAI ; 
 RBJ <= RAJ ; 
 RBK <= RAK ; 
 RBL <= RAL ; 
 RCI <= RBI ; 
 RCJ <= RBJ ; 
 RCK <= RBK ; 
 RCL <= RBL ; 
 RAI <=  KJI & TFB  |  KKI & tfb  ; 
 RAJ <=  KJJ & TFB  |  KKJ & tfb  ; 
 FLI <= ADI ; 
 FLJ <= ADJ ; 
 FLK <= ADK ; 
 FLL <= ADL ; 
 RAO <=  KJO & TFB  |  KKO & tfb  ; 
 RAP <=  KJP & TFB  |  KKP & tfb  ; 
 RAK <=  KJK & TFB  |  KKK & tfb  ; 
 RAL <=  KJL & TFB  |  KKL & tfb  ; 
 FPI <= AHI ; 
 FPJ <= AHJ ; 
 FPK <= AHK ; 
 FPL <= AHL ; 
 kki <= fpi ; 
 kkj <= fpj ; 
 kkk <= fpk ; 
 kkl <= fpl ; 
 kkm <= fpm ; 
 kkn <= fpn ; 
 kko <= fpo ; 
 kkp <= fpp ; 
 kjm <= flm ; 
 kjn <= fln ; 
 kjo <= flo ; 
 kjp <= flp ; 
 RAM <=  KJM & TFB  |  KKM & tfb  ; 
 RAN <=  KJN & TFB  |  KKN & tfb  ; 
 FPM <= AHM ; 
 FPN <= AHN ; 
 FPO <= AHO ; 
 FPP <= AHP ; 
 kji <= fli ; 
 kjj <= flj ; 
 kjk <= flk ; 
 kjl <= fll ; 
 FLM <= ADM ; 
 FLN <= ADN ; 
 FLO <= ADO ; 
 FLP <= ADP ; 
 RBM <= RAM ; 
 RBN <= RAN ; 
 RBO <= RAO ; 
 RBP <= RAP ; 
 RCM <= RBM ; 
 RCN <= RBN ; 
 RCO <= RBO ; 
 RCP <= RBP ; 
 OGI <= RCI ; 
 OGJ <= RCJ ; 
 OGK <= RCK ; 
 OGL <= RCL ; 
 FBC <=  dbc & EBC  |  DBC & ebc  ; 
 FBI <=  dbi & EBC  |  DBI & ebc  ; 
 qgg <= qfc ; 
 qgh <= qfc ; 
 qgi <= qfc ; 
 qgj <= qfc ; 
 FCB <=  dcb & ECB  |  DCB & ecb  ; 
 FCE <=  dce & ECB  |  DCE & ecb  ; 
 FBD <=  dbd & EBD  |  DBD & ebd  ; 
 FBJ <=  dbj & EBD  |  DBJ & ebd  ; 
 OJC <= QHC ; 
 QHC <= QGI ; 
 FBE <=  dbe & EBE  |  DBE & ebe  ; 
 FBK <=  dbk & EBE  |  DBK & ebe  ; 
 GAA <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAE <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAK <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAC <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAI <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAM <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 FBF <=  dbf & EBF  |  DBF & ebf  ; 
 FBL <=  dbl & EBF  |  DBL & ebf  ; 
 GAG <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAL <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAN <=  DAG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAH <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAJ <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAO <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 FCA <=  ECA  ; 
 FCD <=  eca  ; 
 GAB <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAD <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 GAF <=  DDG & EBG & ECH  |  DBG & ECG  |  DCD  ; 
 QJM <=  FLP & fpp  |  flp & FPP  ; 
 OHA <= QJM ; 
 OGM <= RCM ; 
 OGN <= RCN ; 
 OGO <= RCO ; 
 OGP <= RCP ; 
 FCC <=  dcc & ECC  |  DCC & ecc  ; 
 FCF <=  dcf & ECC  |  DCF & ecc  ; 
 BBI <=  IDI  |  ihi & TDF  |  adi & tdf  ; 
 BAI <=  IDI  |  ihi & TDF  |  adi & tdf  ; 
 cai <=  idi  |  IHI & TDF  |  ADI & tdf  ; 
 ADI <=  IDI & TAA  |  IHI & TDA  |  ADI & TCA  ; 
 ADJ <=  IDJ & TAA  |  IHJ & TDA  |  ADJ & TCA  ; 
 BAJ <=  IDJ  |  ihj & TDF  |  adj & tdf  ; 
 caj <=  idj  |  IHJ & TDF  |  ADJ & tdf  ; 
 ahi <= idi ; 
 ahj <= idj ; 
 ahk <= idk ; 
 ahl <= idl ; 
 BAO <=  IDO & jeb  |  iho & TDF  |  ado & tdf  ; 
 cao <=  ido & jeb  |  IHO & TDF  |  ADO & tdf  ; 
 BAK <=  IDK  |  ihk & TDF  |  adk & tdf  ; 
 cak <=  idk  |  IHK & TDF  |  ADK & tdf  ; 
 ADK <=  IDK & TAB  |  IHK & TDB  |  ADK & TCB  ; 
 ADL <=  IDL & TAB  |  IHL & TDB  |  ADL & TCB  ; 
 BAL <=  IDL  |  ihl & TDF  |  adl & tdf  ; 
 cal <=  idl  |  IHL & TDF  |  ADL & tdf  ; 
 ADM <=  IDM & TAC  |  IHM & TDC  |  ADM & TCC  ; 
 ADN <=  IDN & TAC  |  IHN & TDC  |  ADN & TCC  ; 
 BAM <=  IDM  |  ihm & TDF  |  adm & tdf  ; 
 cam <=  idm  |  IHM & TDF  |  ADM & tdf  ; 
 ahm <= idm ; 
 ahn <= idn ; 
 aho <= ido ; 
 BAN <=  IDN  |  ihn & TDF  |  adn & tdf  ; 
 can <=  idn  |  IHN & TDF  |  ADN & tdf  ; 
 ADO <=  IDO & TAD  |  IHO & TDD  |  ADO & TCD  |  TEA  ; 
 DCB <=  CAM  ; 
 DCC <=  CAM  ; 
 BBG <=  IDG  |  ihg & TDH  |  adg & tdh  ; 
 cbg <=  idg  |  IHG & TDH  |  ADG & tdh  ; 
 ADP <=  IDP & TAD  |  IHP & TDD  |  ADP & TCD  ; 
 qja <=  ahp & adp  |  AHP & ADP  ; 
 BBH <=  IDH  |  ihh & TDH  |  adh & tdh  ; 
 cbh <=  idh  |  IHH & TDH  |  ADH & tdh  ; 
 TDA <= QEA & qeb ; 
 TDB <= QEA & qeb ; 
 TDC <= QEA & qeb ; 
 TDD <= QEA & qeb ; 
 ahp <=  idp & tba  |  IDP & TBA  ; 
 RBA <= RAA ; 
 RBB <= RAB ; 
 RBC <= RAC ; 
 RBD <= RAD ; 
 RCA <= RBA ; 
 RCB <= RBB ; 
 RCC <= RBC ; 
 RCD <= RBD ; 
 qfb <= qef & qej ; 
 RAA <=  KJA & TFA  |  KKA & tfa  ; 
 RAB <=  KJB & TFA  |  KKB & tfa  ; 
 QEC <= QDC ; 
 QEF <= QDF ; 
 QEG <= QDG ; 
 QEH <= QDH ; 
 kja <= fla ; 
 kjb <= flb ; 
 kjc <= flc ; 
 kjd <= fld ; 
 RAC <=  KJC & TFA  |  KKC & tfa  ; 
 RAD <=  KJD & TFA  |  KKD & tfa  ; 
 FLA <= ADA ; 
 FLB <= ADB ; 
 FLC <= ADC ; 
 FLD <= ADD ; 
 kka <= fpa ; 
 kkb <= fpb ; 
 kkc <= fpc ; 
 kkd <= fpd ; 
 qfc <= qeg & qek ; 
 FPA <= AHA ; 
 FPB <= AHB ; 
 FPC <= AHC ; 
 FPD <= AHD ; 
 kke <= fpe ; 
 kkf <= fpf ; 
 kkg <= fpg ; 
 kkh <= fph ; 
 QGA <= QFA ; 
 QGB <= QFB ; 
 FPE <= AHE ; 
 FPF <= AHF ; 
 FPG <= AHG ; 
 FPH <= AHH ; 
 kje <= fle ; 
 kjf <= flf ; 
 kjg <= flg ; 
 kjh <= flh ; 
 RAE <=  KJE & TFA  |  KKE & tfa  ; 
 RAF <=  KJF & TFA  |  KKF & tfa  ; 
 FLE <= ADE ; 
 FLF <= ADF ; 
 FLG <= ADG ; 
 FLH <= ADH ; 
 qfa <= qee & qei ; 
 RAG <=  KJG & TFA  |  KKG & tfa  ; 
 RAH <=  KJH & TFA  |  KKH & tfa  ; 
 QEA <= QDA ; 
 QEB <= QDB ; 
 QED <= QDD ; 
 QEE <= QDE ; 
 tba <= qeh & qdh ; 
 RBE <= RAE ; 
 RBF <= RAF ; 
 RBG <= RAG ; 
 RBH <= RAH ; 
 RCE <= RBE ; 
 RCF <= RBF ; 
 RCG <= RBG ; 
 RCH <= RBH ; 
 OGA <= RCA ; 
 OGB <= RCB ; 
 OGC <= RCC ; 
 OGD <= RCD ; 
 FAA <=  EAA  ; 
 FAG <=  eaa  ; 
 FBA <=  EBA  ; 
 FBG <=  eba  ; 
 FAB <=  dab & EAB  |  DAB & eab  ; 
 FAH <=  dah & EAB  |  DAH & eab  ; 
 QYA <= QGB & GAP ; 
 OIA <= QGB & QYA ; 
 gca <=  ZZO & dcd & dag & dbg  |  ZZI & dcd & dag & dbg  |  eag & dag & dbg  |  ebg & dbg & dbg  ; 
 gap <=  ZZO & dag & dbg & dcd  |  ZZI & dag & dbg & dcd  |  ebg & dbg & dcd  |  ecg & dcd & dcd  ; 
 FAE <= dae & EAE |  DAE & eae ; 
 FAK <= dak & EAE |  DAK & eae ; 
 FAD <=  dad & EAD  |  DAD & ead  ; 
 gba <=  ZZO & dbg & dcd & ddg  |  ZZI & dbg & dcd & ddg  |  ech & dcd & ddg  |  eag & ddg & ddg  ; 
 gaq <=  ZZO & ddg & dbg & dcd  |  ZZI & ddg & dbg & dcd  |  ebg & dbg & dcd  |  ecg & dcd & dcd  ; 
 FAF <= daf & EAF |  DAF & eaf ; 
 FAL <= dal & EAF |  DAL & eaf ; 
 OJA <= QHA ; 
 OJB <= QHB ; 
 QHA <= QGA ; 
 QHB <= QGB ; 
 BBC <=  IDC  |  ihc & TDG  |  adc & tdg  ; 
 FAC <=  dac & EAC  |  DAC & eac  ; 
 FAI <=  dai & EAC  |  DAI & eac  ; 
 QEI <= QEA ; 
 QEJ <= QEC ; 
 QEK <= QED ; 
 FAJ <=  daj & EAD  |  DAJ & ead  ; 
 OGE <= RCE ; 
 OGF <= RCF ; 
 OGG <= RCG ; 
 OGH <= RCH ; 
 FBB <=  dbb & EBB  |  DBB & ebb  ; 
 FBH <=  dbh & EBB  |  DBH & ebb  ; 
 BBA <=  IDA  |  iha & TDG  |  ada & tdg  ; 
 cba <=  ida  |  IHA & TDG  |  ADA & tdg  ; 
 BAA <=  IDA  |  iha & TDE  |  ada & tde  ; 
 caa <=  ida  |  IHA & TDE  |  ADA & tde  ; 
 ADA <=  IDA & TAA  |  IHA & TDA  |  ADA & TCA  ; 
 ADB <=  IDB & TAA  |  IHB & TDA  |  ADB & TCA  ; 
 BBB <=  IDB  |  ihb & TDG  |  adb & tdg  ; 
 cbb <=  idb  |  IHB & TDG  |  ADB & tdg  ; 
 BAB <=  IDB  |  ihb & TDE  |  adb & tde  ; 
 cab <=  idb  |  IHB & TDE  |  ADB & tde  ; 
 aha <= ida ; 
 ahb <= idb ; 
 ahc <= idc ; 
 ahd <= idd ; 
 cag <=  idg  |  IHG & TDE  |  ADG & tde  ; 
 BAC <=  IDC  |  ihc & TDE  |  adc & tde  ; 
 cac <=  idc  |  IHC & TDE  |  ADC & tde  ; 
 ADC <=  IDC & TAB  |  IHC & TDB  |  ADC & TCB  ; 
 ADD <=  IDD & TAB  |  IHD & TDB  |  ADD & TCB  ; 
 BAD <=  IDD  |  ihd & TDE  |  add & tde  ; 
 cad <=  idd  |  IHD & TDE  |  ADD & tde  ; 
 ADE <=  IDE & TAC  |  IHE & TDC  |  ADE & TCC  |  TEA  ; 
 BAE <=  IDE  |  ihe & TDE  |  ade & tde  ; 
 cae <=  ide  |  IHE & TDE  |  ADE & tde  ; 
 ADF <=  IDF & TAC  |  IHF & TDC  |  ADF & TCC  |  TEA  ; 
 BAF <=  IDF  |  ihf & TDE  |  adf & tde  ; 
 caf <=  idf  |  IHF & TDE  |  ADF & tde  ; 
 ahe <= ide ; 
 ahf <= idf ; 
 ahg <= idg ; 
 ahh <= idh ; 
 BAG <=  IDG  |  ihg & TDE  |  adg & tde  ; 
 ADG <=  IDG & TAD  |  IHG & TDD  |  ADG & TCD  ; 
 ADH <=  IDH & TAD  |  IHH & TDD  |  ADH & TCD  ; 
 BAH <=  IDH  |  ihh & TDE  |  adh & tde  ; 
 cah <=  idh  |  IHH & TDE  |  ADH & tde  ; 
 TDE <= QEA & qeb ; 
 TDF <= QEA & qeb ; 
 TDG <= QEA & qeb ; 
 TDH <= QEA & qeb ; 
 FKI <= ACI ; 
 FKK <= ACK ; 
 FKL <= ACL ; 
 FKJ <= ACJ ; 
 kfi <=  fki & THA  |  foi & tha  ; 
 kfj <=  fkj & THA  |  foj & tha  ; 
 kfk <=  fkk & THB  |  fok & thb  ; 
 kfl <=  fkl & THB  |  fol & thb  ; 
 FOI <= AGI ; 
 FOJ <= AGJ ; 
 FOK <= AGK ; 
 FOL <= AGL ; 
 kfm <=  fkm & THC  |  fom & thc  ; 
 kfn <=  fkn & THC  |  fon & thc  ; 
 FOM <= AGM ; 
 FON <= AGN ; 
 FOO <= AGO ; 
 FOP <= AGP ; 
 kfo <=  fko & THD  |  foo & thd  ; 
 kfp <=  fkp & THD  |  fop & thd  ; 
 FKM <= ACM ; 
 FKN <= ACN ; 
 FKO <= ACO ; 
 FKP <= ACP ; 
 KCI <=  tuk & tvk & HCI  ; 
 KOI <=  tuk & tvk & HCI  ; 
 KPI <=  tuk & tvk & HCI  ; 
 ofi <=  KFI & TGF  |  kfi & tgf  ; 
 ofj <=  KFJ & TGF  |  kfj & tgf  ; 
 KCJ <=  tuk & tvk & HCJ  ; 
 KOJ <=  tuk & tvk & HCJ  ; 
 KPJ <=  tuk & tvk & HCJ  ; 
 TFA <=  QGH  |  gap  ; 
 TFB <=  QGH  |  gap  ; 
 KCK <=  tuk & tvk & HCK  ; 
 KOK <=  tuk & tvk & HCK  ; 
 KPK <=  tuk & tvk & HCK  ; 
 ofk <=  KFK & TGF  |  kfk & tgf  ; 
 ofl <=  KFL & TGF  |  kfl & tgf  ; 
 KCL <=  tuk & tvk & HCL  ; 
 KOL <=  tuk & tvk & HCL  ; 
 KPL <=  tuk & tvk & HCL  ; 
 KCM <=  tul & tvl & HCM  ; 
 KOM <=  tul & tvl & HCM  ; 
 KPM <=  tul & tvl & HCM  ; 
 ofm <=  KFM & TGF  |  kfm & tgf  ; 
 ofn <=  KFN & TGF  |  kfn & tgf  ; 
 KCN <=  tul & tvl & HCN  ; 
 KON <=  tul & tvl & HCN  ; 
 cbc <=  idc  |  IHC & TDG  |  ADC & tdg  ; 
 KCO <=  tul & tvl & HCO  ; 
 KOO <=  tul & tvl & HCO  ; 
 ofo <=  KFO & TGF  |  kfo & tgf  ; 
 ofp <=  KFP & TGF  |  kfp & tgf  ; 
 KCP <=  tul & tvl & HCP  ; 
 KOP <=  tul & tvl & HCP  ; 
 TOF <= JAB & jba ; 
 TPF <= JAB & JBA ; 
 oci <=  TMF & lfi  |  TNF & lfj  |  TOF & lck  |  TPF & lcl  |  JDB  ; 
 oka <= qkl ; 
 qkj <= qki ; 
 qkk <= qkj ; 
 qkl <= qkk ; 
 TMF <= jab & jaa ; 
 TNF <= jab & JAA ; 
 ocj <=  TMF & lfj  |  TNF & lck  |  TOF & lcl  |  TPF & lcm  |  JDB  ; 
 ocn <=  TMF & lcn  |  TNF & lco  |  TOF & lcp  |  TPF  |  JDA  ; 
 TQK <= jad & jac ; 
 TQL <= jad & jac ; 
 TRK <= jad & JAC ; 
 TRL <= jad & JAC ; 
 ock <=  TMF & lck  |  TNF & lfl  |  TOF & lcm  |  TPF & lcn  |  JDB  ; 
 agi <= ici ; 
 agj <= icj ; 
 agk <= ick ; 
 agl <= icl ; 
 ocl <=  TMF & lfl  |  TNF & lcm  |  TOF & lcn  |  TPF & lco  |  JDB  ; 
 ACK <=  ICK & TAB  |  IGK & TDB  |  ACK & TCB  ; 
 ACL <=  ICL & TAB  |  IGL & TDB  |  ACL & TCB  ; 
 ocm <=  TMF & lcm  |  TNF & lcn  |  TOF & lco  |  TPF & lcp  |  JDA  ; 
 ACM <=  ICM & TAC  |  IGM & TDC  |  ACM & TCC  ; 
 ACN <=  ICN & TAC  |  IGN & TDC  |  ACN & TCC  ; 
 TSK <= JAD & jfc ; 
 TSL <= JAD & jfc ; 
 TTK <= JAD & JFC ; 
 TTL <= JAD & JFC ; 
 agm <= icm ; 
 agn <= icn ; 
 ago <= ico ; 
 agp <= icp ; 
 qkf <= qke ; 
 qkg <= qkf ; 
 qkh <= qkg ; 
 qki <= qkh ; 
 oco <=  TMF & lco  |  TNF & lfp  |  TOF  |  TPF  |  JDA  ; 
 ACO <=  ICO & TAD  |  IGO & TDD  |  ACO & TCD  ; 
 ACP <=  ICP & TAD  |  IGP & TDD  |  ACP & TCD  ; 
 ACI <=  ICI & TAA  |  IGI & TDA  |  ACI & TCA  ; 
 ACJ <=  ICJ & TAA  |  IGJ & TDA  |  ACJ & TCA  ; 
 ocp <=  TMF & lfp  |  TNF  |  TOF  |  TPF  |  JDA  ; 
 TEA <=  QCF  |  QCG  |  QDC  |  QDD  |  JEA  ; 
 FKA <= ACA ; 
 FKB <= ACB ; 
 FKC <= ACC ; 
 FKD <= ACD ; 
 kfb <=  fkb & THA  |  fob & tha  ; 
 kfc <=  fkc & THB  |  foc & thb  ; 
 kfd <=  fkd & THB  |  fod & thb  ; 
 FOA <= AGA ; 
 FOB <= AGB ; 
 FOC <= AGC ; 
 FOD <= AGD ; 
 kfe <=  fke & THC  |  foe & thc  ; 
 kff <=  fkf & THC  |  fof & thc  ; 
 FOE <= AGE ; 
 FOF <= AGF ; 
 FOG <= AGG ; 
 FOH <= AGH ; 
 kfg <=  fkg & THD  |  fog & thd  ; 
 kfh <=  fkh & THD  |  foh & thd  ; 
 kfa <=  fka & THA  |  foa & tha  ; 
 FKE <= ACE ; 
 FKF <= ACF ; 
 FKG <= ACG ; 
 FKH <= ACH ; 
 KCA <=  tui & tvi & HCA  ; 
 KOA <=  tui & tvi & HCA  ; 
 KPA <=  tui & tvi & HCA  ; 
 qbe <=  qab & qab  |  QAD & QAD  ; 
 qbh <=  qad & qab  |  qaa & QAD  |  qac & qaa  ; 
 ofa <=  KFA & TGE  |  kfa & tge  ; 
 ofb <=  KFB & TGE  |  kfb & tge  ; 
 KCB <=  tui & tvi & HCB  ; 
 KOB <=  tui & tvi & HCB  ; 
 KPB <=  tui & tvi & HCB  ; 
 qbf <=  qab  |  qad  |  QAC  ; 
 qbg <=  qab  |  qad  |  qac  ; 
 KCC <=  tui & tvi & HCC  ; 
 KOC <=  tui & tvi & HCC  ; 
 KPC <=  tui & tvi & HCC  ; 
 QXJ <= TVJ & TUJ ; 
 QXK <= TVJ & TUJ ; 
 QXL <= TVJ & TUJ ; 
 ofc <=  KFC & TGE  |  kfc & tge  ; 
 ofd <=  KFD & TGE  |  kfd & tge  ; 
 KCD <=  tui & tvi & HCD  ; 
 KOD <=  tui & tvi & HCD  ; 
 KPD <=  tui & tvi & HCD  ; 
 qxa <=  nca & nba & ncb  ; 
 qxb <=  nca & nba & ncb  ; 
 qxc <=  nca & nba & ncb  ; 
 KCE <=  tuj & tvj & HCE  ; 
 KOE <=  tuj & tvj & HCE  ; 
 KPE <=  tuj & tvj & HCE  ; 
 qba <=  qaa  |  QAE  ; 
 qbb <=  qaa  |  QAE  |  QAC  ; 
 ofe <=  KFE & TGE  |  kfe & tge  ; 
 off <=  KFF & TGE  |  kff & tge  ; 
 KCF <=  tuj & tvj & HCF  ; 
 KOF <=  tuj & tvj & HCF  ; 
 qbc <=  qaa  |  qae  |  QAC  ; 
 qbd <=  qaa  |  gae  |  qac  ; 
 KCG <=  tuj & tvj & HCG  ; 
 KOG <=  tuj & tvj & HCG  ; 
 ofg <=  KFG & TGE  |  kfg & tge  ; 
 ofh <=  KFH & TGE  |  kfh & tge  ; 
 KCH <=  tuj & tvj & HCH  ; 
 KOH <=  tuj & tvj & HCH  ; 
 TOE <= JAB & jba ; 
 TPE <= JAB & JBA ; 
 oca <=  TME & lfa  |  TNE & lfb  |  TOE & lcc  |  TPE & lcd  |  JDD  ; 
 qac <= ijc ; 
 qad <= ijd ; 
 qae <= ije ; 
 TME <= jab & jaa ; 
 TNE <= jab & JAA ; 
 ocb <=  TME & lfb  |  TNE & lcc  |  TOE & lcd  |  TPE & lce  |  JDD  ; 
 ACA <=  ICA & TAA  |  IGA & TDA  |  ACA & TCA  ; 
 ACB <=  ICB & TAA  |  IGB & TDA  |  ACB & TCA  ; 
 TQI <= jad & jac ; 
 TQJ <= jad & jac ; 
 TRI <= jad & JAC ; 
 TRJ <= jad & JAC ; 
 ocg <=  TME & lcg  |  TNE & lfh  |  TOE & lci  |  TPE & lcj  |  JDC  ; 
 occ <=  TME & lcc  |  TNE & lfd  |  TOE & lce  |  TPE & lcf  |  JDD  ; 
 aga <= ica ; 
 agb <= icb ; 
 agc <= icc ; 
 agd <= icd ; 
 ocd <=  TME & lfd  |  TNE & lce  |  TOE & lcf  |  TPE & lcg  |  JDD  ; 
 ACC <=  ICC & TAB  |  IGC & TDB  |  ACC & TCB  ; 
 ACD <=  ICD & TAB  |  IGD & TDB  |  ACD & TCB  ; 
 oce <=  TME & lce  |  TNE & lcf  |  TOE & lcg  |  TPE & lch  |  JDC  ; 
 ACE <=  ICE & TAC  |  IGE & TDC  |  ACE & TCC  ; 
 ACF <=  ICF & TAC  |  IGF & TDC  |  ACF & TCC  ; 
 TSI <= JAD & jfc ; 
 TSJ <= JAD & jfc ; 
 TTI <= JAD & JFC ; 
 TTJ <= JAD & JFC ; 
 ocf <=  TME & lcf  |  TNE & lcg  |  TOE & lch  |  TPE & lci  |  JDC  ; 
 age <= ice ; 
 agf <= icf ; 
 agg <= icg ; 
 agh <= ich ; 
 ACG <=  ICG & TAD  |  IGG & TDD  |  ACG & TCD  ; 
 ACH <=  ICH & TAD  |  IGH & TDD  |  ACH & TCD  ; 
 tge <= qja ; 
 tgf <= qja ; 
 och <=  TME & lfh  |  TNE & lii  |  TOE & lcj  |  TPE & lfk  |  JDC  ; 
 qaa <= ija ; 
 qab <= ijb ; 
 FJI <= ABI ; 
 FJJ <= ABJ ; 
 FJL <= ABL ; 
 FJK <= ABK ; 
 kei <=  fji & THA  |  fni & tha  ; 
 kek <=  fjk & THB  |  fnk & thb  ; 
 kel <=  fjl & THB  |  fnl & thb  ; 
 FNI <= AFI ; 
 FNJ <= AFJ ; 
 FNK <= AFK ; 
 FNL <= AFL ; 
 FJN <= ABN ; 
 FJP <= ABP ; 
 kem <=  fjm & THC  |  fnm & thc  ; 
 ken <=  fjn & THC  |  fnn & thc  ; 
 FNM <= AFM ; 
 FNN <= AFN ; 
 FNO <= AFO ; 
 FNP <= AFP ; 
 keo <=  fjo & THD  |  fno & thd  ; 
 kep <=  fjp & THD  |  fnp & thd  ; 
 kej <=  fjj & THA  |  fnj & tha  ; 
 FJM <= ABM ; 
 FJO <= ABO ; 
 KBI <=  tug & tvg & HBI  |  HCI & TUG  ; 
 KMI <=  tug & tvg & HBI  |  HCI & TUG  ; 
 KNI <=  tug & tvg & HBI  |  HCI & TUG  ; 
 oei <=  KEE & TGD  |  kei & tgd  ; 
 oej <=  KEJ & TGD  |  kej & tgd  ; 
 KBJ <=  tug & tvg & HBJ  |  HCJ & TUG  ; 
 KMJ <=  tug & tvg & HBJ  |  HCJ & TUG  ; 
 KNJ <=  tug & tvg & HBJ  |  HCJ & TUG  ; 
 KBK <=  tug & tvg & HBK  |  HCK & TUG  ; 
 KMK <=  tug & tvg & HBK  |  HCK & TUG  ; 
 KNK <=  tug & tvg & HBK  |  HCK & TUG  ; 
 qxd <=  nbb & nbc & ncc  ; 
 qxe <=  nbb & nbc & ncc  ; 
 qxf <=  nbb & nbc & ncc  ; 
 oek <=  KEK & TGD  |  kek & tgd  ; 
 oel <=  KEL & TGD  |  kel & tgd  ; 
 KBL <=  tug & tvg & HBL  |  HCL & TUG  ; 
 KML <=  tug & tvg & HBL  |  HCL & TUG  ; 
 KNL <=  tug & tvg & HBL  |  HCL & TUG  ; 
 KBM <=  tuh & tvh & HBM  |  HCM & TUH  ; 
 KMM <=  tuh & tvh & HBM  |  HCM & TUH  ; 
 KNM <=  tuh & tvh & HBM  |  HCM & TUH  ; 
 oem <=  KEM & TGD  |  kem & tgd  ; 
 oen <=  KEN & TGD  |  ken & tgd  ; 
 KBN <=  tuh & tvh & HBN  |  HCN & TUH  ; 
 KMN <=  tuh & tvh & HBN  |  HCN & TUH  ; 
 KBO <=  tuh & tvh & HBO  |  HCO & TUH  ; 
 KMO <=  tuh & tvh & HBO  |  HCO & TUH  ; 
 HBK <=  FNK & gag  |  FJK & GAG  ; 
 oeo <=  KEO & TGD  |  keo & tgd  ; 
 oep <=  KEP & TGD  |  kep & tgd  ; 
 KBP <=  tuh & tvh & HBP  |  HCP & TUH  ; 
 KMP <=  tuh & tvh & HBP  |  HCP & TUH  ; 
 TOD <= JAB & jba ; 
 TPD <= JAB & JBA ; 
 obi <=  TMD & lei  |  TND & lej  |  TOD & lbk  |  TPD & lbl  |  JDF  ; 
 TMD <= jab & jaa ; 
 TND <= jab & JAA ; 
 obj <=  TMD & lej  |  TND & lbk  |  TOD & lbl  |  TPD & lbm  |  JDF  ; 
 ABI <=  IBI & TAA  |  IFI & TDA  |  ABI & TCA  ; 
 ABJ <=  IBJ & TAA  |  IFJ & TDA  |  ABJ & TCA  ; 
 TQG <= jbd & jcc ; 
 TQH <= jbd & jbc ; 
 TRG <= jbd & JCC ; 
 TRH <= jbd & JBC ; 
 obk <=  TMD & lbk  |  TND & lel  |  TOD & lbm  |  TPD & lbn  |  JDF  ; 
 afi <= ibi ; 
 afj <= ibj ; 
 afk <= ibk ; 
 afl <= ibl ; 
 obl <=  TMD & lel  |  TND & lbm  |  TOD & lbn  |  TPD & lbo  |  JDF  ; 
 ABK <=  IBK & TAB  |  IFK & TDB  |  ABK & TCB  ; 
 ABL <=  IBL & TAB  |  IFL & TDB  |  ABL & TCB  ; 
 obm <=  TMD & lbm  |  TND & lbn  |  TOD & lbo  |  TPD & lbp  |  JDE  ; 
 ABM <=  IBM & TAC  |  IFM & TDC  |  ABM & TCC  ; 
 ABN <=  IBN & TAC  |  IFN & TDC  |  ABN & TCC  ; 
 TSG <= JBD & jhc ; 
 TSH <= JBD & jgc ; 
 TTG <= JBD & JHC ; 
 TTH <= JBD & JGC ; 
 obn <=  TMD & lbn  |  TND & lbo  |  TOD & lbp  |  TPD & lca  |  JDE  ; 
 afm <= ibm ; 
 afn <= ibn ; 
 afo <= ibo ; 
 afp <= ibp ; 
 qka <= ila ; 
 qkd <= qkc ; 
 qke <= qkd ; 
 obo <=  TMD & lbo  |  TND & lep  |  TOD & lca  |  TPD & lcb  |  JDE  ; 
 ABO <=  IBO & TAD  |  IFO & TDD  |  ABO & TCD  ; 
 ABP <=  IBP & TAD  |  IFP & TDD  |  ABP & TCD  ; 
 qkb <=  qka & QKB  ; 
 QKC <=  QIB & QKB  |  QDI & QKC  ; 
 obp <=  TMD & lep  |  TND & lia  |  TOD & lcb  |  TPD & lfc  |  JDE  ; 
 QIA <=  QAA  |  QAB  ; 
 QIB <=  QIA  ; 
 FJA <= ABA ; 
 FJB <= ABB ; 
 FJC <= ABC ; 
 FJD <= ABD ; 
 kea <=  fja & THE  |  fna & the  ; 
 keb <=  fjb & THE  |  fnb & the  ; 
 kec <=  fjc & THF  |  fnc & thf  ; 
 ked <=  fjd & THF  |  fnd & thf  ; 
 FNA <= AFA ; 
 FNB <= AFB ; 
 FNC <= AFC ; 
 FND <= AFD ; 
 kee <=  fje & THG  |  fne & thg  ; 
 kef <=  fjf & THG  |  fnf & thg  ; 
 FNE <= AFE ; 
 FNF <= AFF ; 
 FNG <= AFG ; 
 FNH <= AFH ; 
 keg <=  fjg & THH  |  fng & thh  ; 
 keh <=  fjh & THH  |  fnh & thh  ; 
 FJE <= ABE ; 
 FJF <= ABF ; 
 FJG <= ABG ; 
 FJH <= ABH ; 
 KBA <=  tue & tve & HBA  |  HCA & TUE  ; 
 KMA <=  tue & tve & HBA  |  HCA & TUE  ; 
 KNA <=  tue & tve & HBA  |  HCA & TUE  ; 
 oea <=  KEA & TGC  |  kea & tgc  ; 
 oeb <=  KEB & TGC  |  keb & tgc  ; 
 KBB <=  tue & tve & HBB  |  HCB & TUE  ; 
 KMB <=  tue & tve & HBB  |  HCB & TUE  ; 
 KNB <=  tue & tve & HBB  |  HCB & TUE  ; 
 oee <=  KEE & TGC  |  kee & tgc  ; 
 KBC <=  tue & tve & HBC  |  HCC & TUE  ; 
 KMC <=  tue & tve & HBC  |  HCC & TUE  ; 
 KNC <=  tue & tve & HBC  |  HCC & TUE  ; 
 qxm <=  qgb & qgc  ; 
 oec <=  KEC & TGC  |  kec & tgc  ; 
 oed <=  KED & TGC  |  ked & tgc  ; 
 KBD <=  tue & tve & HBD  |  HCD & TUE  ; 
 KMD <=  tue & tve & HBD  |  HCD & TUE  ; 
 KND <=  tue & tve & HBD  |  HCD & TUE  ; 
 KBE <=  tuf & tvf & HBE  |  HCE & TUF  ; 
 KME <=  tuf & tvf & HBE  |  HCE & TUF  ; 
 KNE <=  tuf & tvf & HBE  |  HCE & TUF  ; 
 oef <=  KEF & TGC  |  kef & tgc  ; 
 KBF <=  tuf & tvf & HBF  |  HCF & TUF  ; 
 KMF <=  tuf & tvf & HBF  |  HCF & TUF  ; 
 KBG <=  tuf & tvf & HBG  |  HCG & TUF  ; 
 KMG <=  tuf & tvf & HBG  |  HCG & TUF  ; 
 oeg <=  KEG & TGC  |  keg & tgc  ; 
 oeh <=  KEH & TGC  |  keh & tgc  ; 
 KBH <=  tuf & tvf & HBH  |  HCH & TUF  ; 
 KMH <=  tuf & tvf & HBH  |  HCH & TUF  ; 
 TOC <= JAB & jba ; 
 TPC <= JAB & JBA ; 
 oba <=  TMC & lea  |  TNC & leb  |  TOC & lbc  |  TPC & lbd  |  JDH  ; 
 TMC <= jab & jaa ; 
 TNC <= jab & JAA ; 
 obb <=  TMC & leb  |  TNC & lbc  |  TOC & lbd  |  TPC & lbe  |  JDH  ; 
 ABA <=  IBA & TAA  |  IFA & TDA  |  ABA & TCA  ; 
 ABB <=  IBB & TAA  |  IFB & TDA  |  ABB & TCA  ; 
 TQE <= jbd & jcc ; 
 TQF <= jbd & jbc ; 
 TRE <= jbd & JCC ; 
 TRF <= jbd & JBC ; 
 obc <=  TMC & lbc  |  TNC & led  |  TOC & lbe  |  TPC & lbf  |  JDH  ; 
 afa <= iba ; 
 afb <= ibb ; 
 afc <= ibc ; 
 afd <= ibd ; 
 obd <=  TMC & led  |  TNC & lbe  |  TOC & lbf  |  TPC & lbg  |  JDH  ; 
 ABC <=  IBC & TAB  |  IFC & TDB  |  ABC & TCB  ; 
 ABD <=  IBD & TAB  |  IFD & TDB  |  ABD & TCB  ; 
 obe <=  TMC & lbe  |  TNC & lbf  |  TOC & lbg  |  TPC & lbh  |  JDG  ; 
 ABE <=  IBE & TAC  |  IFE & TDC  |  ABE & TCC  ; 
 ABF <=  IBF & TAC  |  IFF & TDC  |  ABF & TCC  ; 
 TSE <= JBD & jhc ; 
 TSF <= JBD & jgc ; 
 TTE <= JBD & JHC ; 
 TTF <= JBD & JGC ; 
 obf <=  TMC & lbf  |  TNC & lbg  |  TOC & lbh  |  TPC & lbi  |  JDG  ; 
 afe <= ibe ; 
 aff <= ibf ; 
 afg <= ibg ; 
 afh <= ibh ; 
 obg <=  TMC & lbg  |  TNC & leh  |  TOC & lbi  |  TPC & lbj  |  JDG  ; 
 ABG <=  IBG & TAD  |  IFG & TDD  |  ABG & TCD  ; 
 ABH <=  IBH & TAD  |  IFH & TDD  |  ABH & TCD  ; 
 tgc <= qja ; 
 tgd <= qja ; 
 obh <=  TMC & leh  |  TNC & lei  |  TOC & lbj  |  TPC & lek  |  JDG  ; 
 FII <= AAI ; 
 FIJ <= AAJ ; 
 FIK <= AAK ; 
 FIL <= AAL ; 
 kdi <=  fii & THE  |  fmi & the  ; 
 kdj <=  fij & THE  |  fmj & the  ; 
 kdk <=  fik & THF  |  fmk & thf  ; 
 kdl <=  fil & THF  |  fml & thf  ; 
 FMI <= AEI ; 
 FMJ <= AEJ ; 
 FMK <= AEK ; 
 FML <= AEL ; 
 kdm <=  fim & THG  |  fmm & thg  ; 
 kdn <=  fin & THG  |  fmn & thg  ; 
 FMM <= AEM ; 
 FMN <= AEN ; 
 FMO <= AEO ; 
 FMP <= AEP ; 
 kdo <=  fio & THH  |  fmo & thh  ; 
 kdp <=  fip & THH  |  fmp & thh  ; 
 FIM <= AAM ; 
 FIN <= AAN ; 
 FIO <= AAO ; 
 FIP <= AAP ; 
 KAI <=  tuc & tvc & HAI  |  HBI & TUC  |  HCI & TVC  ; 
 KLI <=  tuc & tvc & HAI  |  HBI & TUC  |  HCI & TVC  ; 
 odi <=  KDI & TGB  |  kdi & tgb  ; 
 odj <=  KDJ & TGB  |  kdj & tgb  ; 
 KAJ <=  tuc & tvc & HAJ  |  HBJ & TUC  |  HCJ & TVC  ; 
 KLJ <=  tuc & tvc & HAJ  |  HBJ & TUC  |  HCJ & TVC  ; 
 odo <=  KDO & TGB  |  kdo & tgb  ; 
 KAK <=  tuc & tvc & HAK  |  HBK & TUC  |  HCK & TVG  ; 
 KLK <=  tuc & tvc & HAK  |  HBK & TUC  |  HCK & TVG  ; 
 odn <=  KDN & TGB  |  kdn & tgb  ; 
 odk <=  KDK & TGB  |  kdk & tgb  ; 
 odl <=  KDL & TGB  |  kdl & tgb  ; 
 KAL <=  tuc & tvc & HAL  |  HBL & TUC  |  HCL & TVG  ; 
 KLL <=  tuc & tvc & HAL  |  HBL & TUC  |  HCL & TVG  ; 
 KQL <=  tuc & tvc & HAL  |  HBL & TUC  |  HCL & TVG  ; 
 qxg <=  nbd & nbe & nbf  ; 
 qxh <=  nbd & nbe & nbf  ; 
 qxi <=  nbd & nbe & nbf  ; 
 KAM <=  tud & tvd & HAM  |  HBM & TUD  |  HCM & TVD  ; 
 KLM <=  tud & tvd & HAM  |  HBM & TUD  |  HCM & TVD  ; 
 KQM <=  tud & tvd & HAM  |  HBM & TUD  |  HCM & TVD  ; 
 odm <=  KDM & TGB  |  kdm & tgb  ; 
 KLN <=  tud & tvd & HAN  |  HBN & TUD  |  HCN & TVD  ; 
 KAO <=  tud & tvd & HAO  |  HBO & TUD  |  HCO & TVD  ; 
 KLO <=  tud & tvd & HAO  |  HBO & TUD  |  HCO & TVD  ; 
 KAN <=  tud & tvd & HAN  |  HBN & TUD  |  HCN & TVD  ; 
 odp <=  KDP & TGB  |  kdp & tgb  ; 
 KAP <=  tud & tvd & HAP  |  HBP & TUD  |  HCP & TVD  ; 
 KLP <=  tud & tvd & HAP  |  HBP & TUD  |  HCP & TVD  ; 
 TOB <= JBB & jca ; 
 TPB <= JBB & JCA ; 
 oai <=  TMB & ldi  |  TNB & ldj  |  TOB & lak  |  TPB & lal  |  JDJ  ; 
 oar <=  TMA & lar  |  TNA & laa  |  TOA & lab  |  TPA & ldc  |  JDM  ; 
 TMB <= jbb & jaa ; 
 TNB <= jbb & JAA ; 
 oaj <=  TMB & ldj  |  TNB & lak  |  TOB & lal  |  TPB & lam  |  JDJ  ; 
 AAI <=  IAI & TAA  |  IEI & TDA  |  AAI & TCA  ; 
 AAJ <=  IAJ & TAA  |  IEJ & TDA  |  AAJ & TCA  ; 
 TQC <= jcd & jcc ; 
 TQD <= jcd & jbc ; 
 TRC <= jcd & JCC ; 
 TRD <= jcd & JBC ; 
 oao <=  TMB & ldo  |  TNB & ldp  |  TOB & lba  |  TPB & lbb  |  JDI  ; 
 oak <=  TMB & lak  |  TNB & ldl  |  TOB & lam  |  TPB & lan  |  JDJ  ; 
 aei <= iai ; 
 aej <= iaj ; 
 aek <= iak ; 
 ael <= ial ; 
 QGC <= QFC ; 
 QGD <= QFC ; 
 QGE <= QFC ; 
 QGF <= QFC ; 
 oal <=  TMB & ldl  |  TNB & lam  |  TOB & lan  |  TPB & lao  |  JDJ  ; 
 AAK <=  IAK & TAB  |  IEK & TDB  |  AAK & TCB  ; 
 AAL <=  IAL & TAB  |  IEL & TDB  |  AAL & TCB  ; 
 tqm <=  JHC  |  JCD  ; 
 tqn <=  JHC  |  JCD  ; 
 tqo <=  JHC  |  JCD  ; 
 oam <=  TMB & lam  |  TNB & lan  |  TOB & lao  |  TPB & lap  |  JDI  ; 
 AAM <=  IAM & TAC  |  IEM & TDC  |  AAM & TCC  ; 
 AAN <=  IAN & TAC  |  IEN & TDC  |  AAN & TCC  ; 
 TSC <= JBD & jhc ; 
 TSD <= JBD & jgc ; 
 TTC <= JBD & JHC ; 
 TTD <= JBD & JGC ; 
 oan <=  TMB & lan  |  TNB & ldo  |  TOB & lap  |  TPB & lba  |  JDI  ; 
 aem <= iam ; 
 aen <= ian ; 
 aeo <= iao ; 
 aep <= iap ; 
 kar <=  TVK & TUK & TUK & TVK  |  hap & TUK & TVK  |  hbp & TVK  |  tvd & tud  ; 
 AAP <=  IAP & TAD  |  IEP & TDD  |  AAP & TCD  ; 
 AAO <=  IAO & TAD  |  IEO & TDD  |  AAO & TCD  ; 
 KAQ <=  HCP & TUK & TVK  ; 
 oap <=  TMB & ldp  |  TNB & lha  |  TOB & lbb  |  TPB & lec  |  JDI  ; 
 qdi <= qci ; 
 KAA <=  tua & tva & HAA  |  HBA & TUA  |  HCA & TVA  ; 
 QDC <=  QCC & QCI  |  QDC & QCI  ; 
 QDF <= QCF ; 
 QDG <= QCG ; 
 KAB <=  tua & tva & HAB  |  HBB & TUA  |  HCB & TVA  ; 
 QDD <=  QCD & QCI  |  QDD & QCI  ; 
 kda <=  fia & THE  |  fma & the  ; 
 kdb <=  fib & THE  |  fmb & the  ; 
 FIA <= AAA ; 
 FIB <= AAB ; 
 FIC <= AAC ; 
 FID <= AAD ; 
 KAC <=  tua & tva & HAC  |  HBC & TUA  |  HCC & TVE  ; 
 KAE <=  tub & tvb & HAE  |  HBE & TUI  |  HCE & TVF  ; 
 kdc <=  fic & THF  |  fmc & thf  ; 
 kdd <=  fid & THF  |  fmd & thf  ; 
 FMA <= AEA ; 
 FMB <= AEB ; 
 FMC <= AEC ; 
 FMD <= AED ; 
 KAD <=  tua & tva & HAD  |  HBD & TUA  |  HCD & TVE  ; 
 kde <=  fie & THG  |  fme & thg  ; 
 kdf <=  fif & THG  |  fmf & thg  ; 
 FME <= AEE ; 
 FMF <= AEF ; 
 FMG <= AEG ; 
 FMH <= AEH ; 
 kdg <=  fig & THH  |  fmg & thh  ; 
 kdh <=  fih & THH  |  fmh & thh  ; 
 FIE <= AAE ; 
 FIF <= AAF ; 
 FIG <= AAG ; 
 FIH <= AAH ; 
 QDH <=  QDH & QCI  |  QCH  ; 
 QDA <=  QCA & QCI  |  QDA & QCI  ; 
 QDB <=  QCB & QCI  |  QDB & QCI  ; 
 QCA <= QBA ; 
 QCB <= QBB ; 
 QCD <= QBD ; 
 QCE <= QBE ; 
 QDE <= QCE ; 
 QCI <= IKA ; 
 QCC <= QBC ; 
 QCF <= QBF ; 
 QCG <= QBG ; 
 QCH <= QBH ; 
 oda <=  KDA & TGA  |  kda & tga  ; 
 odb <=  KDB & TGA  |  kdb & tga  ; 
 odc <=  KDC & TGA  |  kdc & tga  ; 
 odd <=  KDD & TGA  |  kdd & tga  ; 
 KLD <=  tua & tva & HAD  |  HBD & TUA  |  HCD & TVE  ; 
 ode <=  KDE & TGA  |  kde & tga  ; 
 odf <=  KDF & TGA  |  kdf & tga  ; 
 KAF <=  tub & tvb & HAF  |  HBF & TUI  |  HCF & TVF  ; 
 qdj <= qdb ; 
 KAG <=  tub & tvb & HAG  |  HBG & TUB  |  HCG & TVB  ; 
 odg <=  KDG & TGA  |  kdg & tga  ; 
 odh <=  KDH & TGA  |  kdh & tga  ; 
 KAH <=  tub & tvb & HAH  |  HBH & TUB  |  HCH & TVB  ; 
 KLH <=  tub & tvb & HAH  |  HBH & TUB  |  HCH & TVB  ; 
 TOA <= JBB & jca ; 
 TPA <= JBB & JCA ; 
 oaa <=  TMA & laa  |  TNA & lab  |  TOA & lac  |  TPA & lad  |  JDL  ; 
 taa <= qce & qcb ; 
 tab <= qce & qcb ; 
 tac <= qce & qcb ; 
 tad <= qce & qcb ; 
 TMA <= jbb & jca ; 
 TNA <= jbb & JCA ; 
 oab <=  TMA & lab  |  TNA & lac  |  TOA & lad  |  TPA & lae  |  JDL  ; 
 AAA <=  IAA & TAA  |  IEA & TDA  |  AAA & TCA  ; 
 AAB <=  IAB & TAA  |  IEB & TDA  |  AAB & TCA  ; 
 TQA <= jcd & jcc ; 
 TQB <= jcd & jbc ; 
 TRA <= jcd & JCC ; 
 TRB <= jcd & JBC ; 
 oag <=  TMA & lag  |  TNA & ldh  |  TOA & lai  |  TPA & laj  |  JDK  ; 
 oac <=  TMA & lac  |  TNA & ldd  |  TOA & lae  |  TPA & laf  |  JDL  ; 
 aea <= iaa ; 
 aeb <= iab ; 
 aec <= iac ; 
 aed <= iad ; 
 oad <=  TMA & ldd  |  TNA & lae  |  TOA & laf  |  TPA & lag  |  JDL  ; 
 AAC <=  IAC & TAB  |  IEC & TDB  |  AAC & TCB  ; 
 AAD <=  IAD & TAB  |  IED & TDB  |  AAD & TCB  ; 
 oae <=  TMA & lae  |  TNA & laf  |  TOA & lag  |  TPA & lah  |  JDK  ; 
 AAE <=  IAE & TAC  |  IEE & TDC  |  AAE & TCC  ; 
 AAF <=  IAF & TAC  |  IEF & TDC  |  AAF & TCC  ; 
 TSA <= JBD & jhc ; 
 TSB <= JBD & jgc ; 
 TTA <= JBD & JHC ; 
 TTB <= JBD & JGC ; 
 oaf <=  TMA & laf  |  TNA & lag  |  TOA & lah  |  TPA & lai  |  JDK  ; 
 aee <= iae ; 
 aef <= iaf ; 
 aeg <= iag ; 
 aeh <= iah ; 
 AAG <=  IAG & TAD  |  IEG & TDD  |  AAG & TCD  ; 
 AAH <=  IAH & TAD  |  IEH & TDD  |  AAH & TCD  ; 
 tga <= qja ; 
 tgb <= qja ; 
 oah <=  TMA & ldh  |  TNA & lgi  |  TOA & laj  |  TPA & ldk  |  JDK  ; 
 tca <= jia & qde ; 
 tcb <= jia & qde ; 
 tcc <= jia & qde ; 
 tcd <= jia & qde ; 
 end 
end module
