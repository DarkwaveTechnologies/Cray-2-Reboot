module eb( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFF, 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IHA, 
 IHB, 
 IHC, 
 IIA, 
 IIB, 
 IJA, 
 IJB, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IKI, 
 IKJ, 
 IKK, 
 IKL, 
 IKM, 
 IKN, 
 IKO, 
 IKP, 
 IKQ, 
 IKR, 
 IKS, 
 IKT, 
 IMA, 
 INA, 
 INB, 
 INC, 
 IND, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OKN, 
 OKO, 
 OKP, 
 OKQ, 
 OKR, 
 OKS, 
 OKT, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
OLH ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFF; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IIA; 
 input IIB; 
 input IJA; 
 input IJB; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IKI; 
 input IKJ; 
 input IKK; 
 input IKL; 
 input IKM; 
 input IKN; 
 input IKO; 
 input IKP; 
 input IKQ; 
 input IKR; 
 input IKS; 
 input IKT; 
 input IMA; 
 input INA; 
 input INB; 
 input INC; 
 input IND; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OKN; 
 output OKO; 
 output OKP; 
 output OKQ; 
 output OKR; 
 output OKS; 
 output OKT; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aae ;
reg  aaf ;
reg  aag ;
reg  aah ;
reg  aai ;
reg  aaj ;
reg  aak ;
reg  aal ;
reg  aam ;
reg  aan ;
reg  aao ;
reg  aap ;
reg  aar ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  abe ;
reg  abf ;
reg  abg ;
reg  abh ;
reg  abi ;
reg  abj ;
reg  abk ;
reg  abl ;
reg  abm ;
reg  abn ;
reg  abo ;
reg  abp ;
reg  baa ;
reg  bab ;
reg  bac ;
reg  bad ;
reg  bae ;
reg  baf ;
reg  bag ;
reg  bah ;
reg  bai ;
reg  baj ;
reg  bak ;
reg  bal ;
reg  bam ;
reg  ban ;
reg  bao ;
reg  bap ;
reg  bba ;
reg  bbb ;
reg  bbc ;
reg  bbd ;
reg  bbe ;
reg  bbf ;
reg  bbg ;
reg  bbh ;
reg  bbi ;
reg  bbj ;
reg  bbk ;
reg  bbl ;
reg  bbm ;
reg  bbn ;
reg  bbo ;
reg  bbp ;
reg  bca ;
reg  bcb ;
reg  bcc ;
reg  bcd ;
reg  bce ;
reg  bcf ;
reg  bcg ;
reg  bch ;
reg  bci ;
reg  bcj ;
reg  bck ;
reg  bcl ;
reg  bcm ;
reg  bcn ;
reg  bco ;
reg  bcp ;
reg  bda ;
reg  bdb ;
reg  bdc ;
reg  bdd ;
reg  bde ;
reg  bdf ;
reg  bdg ;
reg  bdh ;
reg  bdi ;
reg  bdj ;
reg  bdk ;
reg  bdl ;
reg  bdm ;
reg  bdn ;
reg  bdo ;
reg  bdp ;
reg  caj ;
reg  cak ;
reg  cal ;
reg  cam ;
reg  can ;
reg  cao ;
reg  cap ;
reg  cbj ;
reg  cbk ;
reg  cbl ;
reg  cbm ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DDA ;
reg  DDB ;
reg  DDC ;
reg  DDD ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EAI ;
reg  EAJ ;
reg  EAK ;
reg  EAL ;
reg  EAM ;
reg  EAN ;
reg  EAO ;
reg  EAP ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBH ;
reg  EBI ;
reg  EBJ ;
reg  EBK ;
reg  EBL ;
reg  EBM ;
reg  EBN ;
reg  EBO ;
reg  EBP ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GAI ;
reg  GAJ ;
reg  GAK ;
reg  GAL ;
reg  GAM ;
reg  GAN ;
reg  GAO ;
reg  GAP ;
reg  GBA ;
reg  GBB ;
reg  GBC ;
reg  GBD ;
reg  GBE ;
reg  GBF ;
reg  GBG ;
reg  GBH ;
reg  GBI ;
reg  GBJ ;
reg  GBK ;
reg  GBL ;
reg  GBM ;
reg  GBN ;
reg  GBO ;
reg  GBP ;
reg  GCA ;
reg  GCB ;
reg  GCC ;
reg  GCD ;
reg  GCE ;
reg  GCF ;
reg  GCG ;
reg  GCH ;
reg  GCI ;
reg  GCJ ;
reg  GCK ;
reg  GCL ;
reg  GCM ;
reg  GCN ;
reg  GCO ;
reg  GCP ;
reg  GDA ;
reg  GDB ;
reg  GDC ;
reg  GDD ;
reg  GDE ;
reg  GDF ;
reg  GDG ;
reg  GDH ;
reg  GDI ;
reg  GDJ ;
reg  GDK ;
reg  GDL ;
reg  GDM ;
reg  GDN ;
reg  GDO ;
reg  GDP ;
reg  haa ;
reg  hab ;
reg  hac ;
reg  had ;
reg  hae ;
reg  haf ;
reg  hag ;
reg  hah ;
reg  hai ;
reg  haj ;
reg  hak ;
reg  hal ;
reg  ham ;
reg  han ;
reg  hao ;
reg  hap ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hbf ;
reg  hbg ;
reg  hbh ;
reg  hbi ;
reg  hbj ;
reg  hbk ;
reg  hbl ;
reg  hbm ;
reg  hbn ;
reg  hbo ;
reg  hbp ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hce ;
reg  hcf ;
reg  hcg ;
reg  hch ;
reg  hci ;
reg  hcj ;
reg  hck ;
reg  hcl ;
reg  hcm ;
reg  hcn ;
reg  hco ;
reg  hcp ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  hdf ;
reg  hdg ;
reg  hdh ;
reg  hdi ;
reg  hdj ;
reg  hdk ;
reg  hdl ;
reg  hdm ;
reg  hdn ;
reg  hdo ;
reg  hdp ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LAG ;
reg  LAH ;
reg  LAI ;
reg  LAJ ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  LBI ;
reg  LBJ ;
reg  LBK ;
reg  LBL ;
reg  LBM ;
reg  LBN ;
reg  LCA ;
reg  LCB ;
reg  LCC ;
reg  LCD ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  MCA ;
reg  MCB ;
reg  MCC ;
reg  mda ;
reg  mdb ;
reg  mdc ;
reg  mdd ;
reg  MDE ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NCG ;
reg  NCH ;
reg  NCI ;
reg  NCJ ;
reg  NCK ;
reg  NCL ;
reg  NCM ;
reg  NCN ;
reg  NCO ;
reg  NCP ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NDE ;
reg  NDF ;
reg  NDG ;
reg  NDH ;
reg  NDI ;
reg  NDJ ;
reg  NDK ;
reg  NDL ;
reg  NDM ;
reg  NDN ;
reg  NDO ;
reg  NDP ;
reg  oaa ;
reg  oab ;
reg  oac ;
reg  oad ;
reg  oae ;
reg  oaf ;
reg  oag ;
reg  oah ;
reg  oai ;
reg  oaj ;
reg  oak ;
reg  oal ;
reg  oam ;
reg  oan ;
reg  oao ;
reg  oap ;
reg  oba ;
reg  obb ;
reg  obc ;
reg  obd ;
reg  obe ;
reg  obf ;
reg  obg ;
reg  obh ;
reg  obi ;
reg  obj ;
reg  obk ;
reg  obl ;
reg  obm ;
reg  obn ;
reg  obo ;
reg  obp ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  odk ;
reg  odl ;
reg  odm ;
reg  odn ;
reg  odo ;
reg  odp ;
reg  oea ;
reg  oeb ;
reg  oec ;
reg  oed ;
reg  oee ;
reg  oef ;
reg  oeg ;
reg  oeh ;
reg  oei ;
reg  oej ;
reg  oek ;
reg  oel ;
reg  oem ;
reg  oen ;
reg  oeo ;
reg  oep ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  ofe ;
reg  off ;
reg  ofg ;
reg  ofh ;
reg  ofi ;
reg  ofj ;
reg  ofk ;
reg  ofl ;
reg  ofm ;
reg  ofn ;
reg  ofo ;
reg  ofp ;
reg  OGA ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  OKG ;
reg  OKH ;
reg  OKI ;
reg  OKJ ;
reg  OKK ;
reg  OKL ;
reg  OKM ;
reg  OKN ;
reg  OKO ;
reg  OKP ;
reg  okq ;
reg  OKR ;
reg  OKS ;
reg  OKT ;
reg  OLA ;
reg  olb ;
reg  olc ;
reg  old ;
reg  ole ;
reg  OLF ;
reg  OLG ;
reg  olh ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAI ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PAN ;
reg  PAO ;
reg  PAP ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PCO ;
reg  PCP ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PDJ ;
reg  PDK ;
reg  PDL ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  PDP ;
reg  qaa ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  qak ;
reg  qal ;
reg  QAM ;
reg  QAN ;
reg  QAO ;
reg  QAP ;
reg  qaq ;
reg  QAT ;
reg  QBA ;
reg  QBB ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCE ;
reg  QCF ;
reg  QCG ;
reg  QCH ;
reg  QCI ;
reg  QCJ ;
reg  QCK ;
reg  QCL ;
reg  QCM ;
reg  QCN ;
reg  QCO ;
reg  QCP ;
reg  QCQ ;
reg  QCR ;
reg  QCS ;
reg  QCT ;
reg  QCU ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QDF ;
reg  QDG ;
reg  QDH ;
reg  QDI ;
reg  QDJ ;
reg  QDK ;
reg  QDL ;
reg  QDM ;
reg  QDN ;
reg  QDO ;
reg  QEA ;
reg  QEB ;
reg  QFA ;
reg  QFB ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  QGE ;
reg  QGF ;
reg  QHA ;
reg  QHB ;
reg  QHC ;
reg  QHD ;
reg  QHE ;
reg  QIA ;
reg  QIB ;
reg  QJA ;
reg  QJB ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QKD ;
reg  QKE ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  QMA ;
reg  QMB ;
reg  QMC ;
reg  QMD ;
reg  qme ;
reg  QMF ;
reg  QMG ;
reg  qmh ;
reg  QMI ;
reg  QMJ ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  QND ;
reg  qoa ;
reg  qob ;
reg  qoc ;
reg  QOD ;
reg  QPA ;
reg  QPB ;
reg  QPC ;
reg  QPD ;
reg  QPE ;
reg  QPF ;
reg  QPG ;
reg  QPH ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QQD ;
reg  QQE ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  QRF ;
reg  QRG ;
reg  QRH ;
reg  QRI ;
reg  QRJ ;
reg  QRK ;
reg  QRL ;
reg  QRM ;
reg  QRN ;
reg  QRO ;
reg  QRP ;
reg  QSA ;
reg  QSB ;
reg  QSC ;
reg  QSD ;
reg  QSE ;
reg  QSF ;
reg  QSG ;
reg  QSH ;
reg  QSI ;
reg  QSJ ;
reg  QSK ;
reg  QSL ;
reg  QSM ;
reg  QSN ;
reg  QSO ;
reg  QSP ;
reg  QTA ;
reg  QTB ;
reg  QTC ;
reg  QTD ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QUD ;
reg  que ;
reg  quf ;
reg  QUG ;
reg  QUH ;
reg  QVA ;
reg  QVB ;
reg  QVC ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  SAD ;
reg  SAE ;
reg  SAF ;
reg  SAG ;
reg  SAH ;
reg  SAI ;
reg  SAJ ;
reg  SAK ;
reg  SAL ;
reg  uaa ;
reg  uab ;
reg  uac ;
reg  uad ;
reg  uae ;
reg  uaf ;
reg  uag ;
reg  uah ;
reg  uai ;
reg  uaj ;
reg  uak ;
reg  ual ;
reg  uam ;
reg  uan ;
reg  uao ;
reg  uap ;
reg  uba ;
reg  ubb ;
reg  ubc ;
reg  ubd ;
reg  ube ;
reg  ubf ;
reg  ubg ;
reg  ubh ;
reg  ubi ;
reg  ubj ;
reg  ubk ;
reg  ubl ;
reg  ubm ;
reg  ubn ;
reg  ubo ;
reg  ubp ;
reg  uca ;
reg  ucb ;
reg  ucc ;
reg  ucd ;
reg  uce ;
reg  ucf ;
reg  ucg ;
reg  uch ;
reg  uci ;
reg  ucj ;
reg  uck ;
reg  ucl ;
reg  ucm ;
reg  ucn ;
reg  uco ;
reg  ucp ;
reg  uda ;
reg  udb ;
reg  udc ;
reg  udd ;
reg  ude ;
reg  udf ;
reg  udg ;
reg  udh ;
reg  udi ;
reg  udj ;
reg  udk ;
reg  udl ;
reg  udm ;
reg  udn ;
reg  udo ;
reg  udp ;
reg  vaa ;
reg  vab ;
reg  VAC ;
reg  VAD ;
reg  vba ;
reg  vbb ;
reg  VBC ;
reg  VBD ;
reg  vca ;
reg  vcb ;
reg  VCC ;
reg  VCD ;
reg  vda ;
reg  vdb ;
reg  VDC ;
reg  VDD ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WAI ;
reg  WAJ ;
reg  WAK ;
reg  WAL ;
reg  WAM ;
reg  WAN ;
reg  WAO ;
reg  WAP ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WBI ;
reg  WBJ ;
reg  WBK ;
reg  WBL ;
reg  WBM ;
reg  WBN ;
reg  WBO ;
reg  WBP ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WCI ;
reg  WCJ ;
reg  WCK ;
reg  WCL ;
reg  WCM ;
reg  WCN ;
reg  WCO ;
reg  WCP ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WDI ;
reg  WDJ ;
reg  WDK ;
reg  WDL ;
reg  WDM ;
reg  WDN ;
reg  WDO ;
reg  WDP ;
reg  XAA ;
reg  XAB ;
reg  XAC ;
reg  XAD ;
reg  XAE ;
reg  XAF ;
reg  XAG ;
reg  XAH ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  AAE ;
wire  AAF ;
wire  AAG ;
wire  AAH ;
wire  AAI ;
wire  AAJ ;
wire  AAK ;
wire  AAL ;
wire  AAM ;
wire  AAN ;
wire  AAO ;
wire  AAP ;
wire  AAR ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ABE ;
wire  ABF ;
wire  ABG ;
wire  ABH ;
wire  ABI ;
wire  ABJ ;
wire  ABK ;
wire  ABL ;
wire  ABM ;
wire  ABN ;
wire  ABO ;
wire  ABP ;
wire  BAA ;
wire  BAB ;
wire  BAC ;
wire  BAD ;
wire  BAE ;
wire  BAF ;
wire  BAG ;
wire  BAH ;
wire  BAI ;
wire  BAJ ;
wire  BAK ;
wire  BAL ;
wire  BAM ;
wire  BAN ;
wire  BAO ;
wire  BAP ;
wire  BBA ;
wire  BBB ;
wire  BBC ;
wire  BBD ;
wire  BBE ;
wire  BBF ;
wire  BBG ;
wire  BBH ;
wire  BBI ;
wire  BBJ ;
wire  BBK ;
wire  BBL ;
wire  BBM ;
wire  BBN ;
wire  BBO ;
wire  BBP ;
wire  BCA ;
wire  BCB ;
wire  BCC ;
wire  BCD ;
wire  BCE ;
wire  BCF ;
wire  BCG ;
wire  BCH ;
wire  BCI ;
wire  BCJ ;
wire  BCK ;
wire  BCL ;
wire  BCM ;
wire  BCN ;
wire  BCO ;
wire  BCP ;
wire  BDA ;
wire  BDB ;
wire  BDC ;
wire  BDD ;
wire  BDE ;
wire  BDF ;
wire  BDG ;
wire  BDH ;
wire  BDI ;
wire  BDJ ;
wire  BDK ;
wire  BDL ;
wire  BDM ;
wire  BDN ;
wire  BDO ;
wire  BDP ;
wire  CAJ ;
wire  CAK ;
wire  CAL ;
wire  CAM ;
wire  CAN ;
wire  CAO ;
wire  CAP ;
wire  CBJ ;
wire  CBK ;
wire  CBL ;
wire  CBM ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dda ;
wire  ddb ;
wire  ddc ;
wire  ddd ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eai ;
wire  eaj ;
wire  eak ;
wire  eal ;
wire  eam ;
wire  ean ;
wire  eao ;
wire  eap ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebh ;
wire  ebi ;
wire  ebj ;
wire  ebk ;
wire  ebl ;
wire  ebm ;
wire  ebn ;
wire  ebo ;
wire  ebp ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fam ;
wire  FAM ;
wire  fan ;
wire  FAN ;
wire  fao ;
wire  FAO ;
wire  fap ;
wire  FAP ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  fbi ;
wire  FBI ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbl ;
wire  FBL ;
wire  fbm ;
wire  FBM ;
wire  fbn ;
wire  FBN ;
wire  fbo ;
wire  FBO ;
wire  fbp ;
wire  FBP ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fcg ;
wire  FCG ;
wire  fch ;
wire  FCH ;
wire  fci ;
wire  FCI ;
wire  fcj ;
wire  FCJ ;
wire  fck ;
wire  FCK ;
wire  fcl ;
wire  FCL ;
wire  fcm ;
wire  FCM ;
wire  fcn ;
wire  FCN ;
wire  fco ;
wire  FCO ;
wire  fcp ;
wire  FCP ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fdh ;
wire  FDH ;
wire  fdi ;
wire  FDI ;
wire  fdj ;
wire  FDJ ;
wire  fdk ;
wire  FDK ;
wire  fdl ;
wire  FDL ;
wire  fdm ;
wire  FDM ;
wire  fdn ;
wire  FDN ;
wire  fdo ;
wire  FDO ;
wire  fdp ;
wire  FDP ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gai ;
wire  gaj ;
wire  gak ;
wire  gal ;
wire  gam ;
wire  gan ;
wire  gao ;
wire  gap ;
wire  gba ;
wire  gbb ;
wire  gbc ;
wire  gbd ;
wire  gbe ;
wire  gbf ;
wire  gbg ;
wire  gbh ;
wire  gbi ;
wire  gbj ;
wire  gbk ;
wire  gbl ;
wire  gbm ;
wire  gbn ;
wire  gbo ;
wire  gbp ;
wire  gca ;
wire  gcb ;
wire  gcc ;
wire  gcd ;
wire  gce ;
wire  gcf ;
wire  gcg ;
wire  gch ;
wire  gci ;
wire  gcj ;
wire  gck ;
wire  gcl ;
wire  gcm ;
wire  gcn ;
wire  gco ;
wire  gcp ;
wire  gda ;
wire  gdb ;
wire  gdc ;
wire  gdd ;
wire  gde ;
wire  gdf ;
wire  gdg ;
wire  gdh ;
wire  gdi ;
wire  gdj ;
wire  gdk ;
wire  gdl ;
wire  gdm ;
wire  gdn ;
wire  gdo ;
wire  gdp ;
wire  HAA ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  HAE ;
wire  HAF ;
wire  HAG ;
wire  HAH ;
wire  HAI ;
wire  HAJ ;
wire  HAK ;
wire  HAL ;
wire  HAM ;
wire  HAN ;
wire  HAO ;
wire  HAP ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HBF ;
wire  HBG ;
wire  HBH ;
wire  HBI ;
wire  HBJ ;
wire  HBK ;
wire  HBL ;
wire  HBM ;
wire  HBN ;
wire  HBO ;
wire  HBP ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HCE ;
wire  HCF ;
wire  HCG ;
wire  HCH ;
wire  HCI ;
wire  HCJ ;
wire  HCK ;
wire  HCL ;
wire  HCM ;
wire  HCN ;
wire  HCO ;
wire  HCP ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  HDF ;
wire  HDG ;
wire  HDH ;
wire  HDI ;
wire  HDJ ;
wire  HDK ;
wire  HDL ;
wire  HDM ;
wire  HDN ;
wire  HDO ;
wire  HDP ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iff ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  iia ;
wire  iib ;
wire  ija ;
wire  ijb ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  iki ;
wire  ikj ;
wire  ikk ;
wire  ikl ;
wire  ikm ;
wire  ikn ;
wire  iko ;
wire  ikp ;
wire  ikq ;
wire  ikr ;
wire  iks ;
wire  ikt ;
wire  ima ;
wire  ina ;
wire  inb ;
wire  inc ;
wire  ind ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgg ;
wire  JGG ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jja ;
wire  JJA ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jke ;
wire  JKE ;
wire  jkf ;
wire  JKF ;
wire  jkg ;
wire  JKG ;
wire  jkh ;
wire  JKH ;
wire  jki ;
wire  JKI ;
wire  jkj ;
wire  JKJ ;
wire  jkk ;
wire  JKK ;
wire  jkl ;
wire  JKL ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lag ;
wire  lah ;
wire  lai ;
wire  laj ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  lbi ;
wire  lbj ;
wire  lbk ;
wire  lbl ;
wire  lbm ;
wire  lbn ;
wire  lca ;
wire  lcb ;
wire  lcc ;
wire  lcd ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  mca ;
wire  mcb ;
wire  mcc ;
wire  MDA ;
wire  MDB ;
wire  MDC ;
wire  MDD ;
wire  mde ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  ncg ;
wire  nch ;
wire  nci ;
wire  ncj ;
wire  nck ;
wire  ncl ;
wire  ncm ;
wire  ncn ;
wire  nco ;
wire  ncp ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nde ;
wire  ndf ;
wire  ndg ;
wire  ndh ;
wire  ndi ;
wire  ndj ;
wire  ndk ;
wire  ndl ;
wire  ndm ;
wire  ndn ;
wire  ndo ;
wire  ndp ;
wire  OAA ;
wire  OAB ;
wire  OAC ;
wire  OAD ;
wire  OAE ;
wire  OAF ;
wire  OAG ;
wire  OAH ;
wire  OAI ;
wire  OAJ ;
wire  OAK ;
wire  OAL ;
wire  OAM ;
wire  OAN ;
wire  OAO ;
wire  OAP ;
wire  OBA ;
wire  OBB ;
wire  OBC ;
wire  OBD ;
wire  OBE ;
wire  OBF ;
wire  OBG ;
wire  OBH ;
wire  OBI ;
wire  OBJ ;
wire  OBK ;
wire  OBL ;
wire  OBM ;
wire  OBN ;
wire  OBO ;
wire  OBP ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  ODK ;
wire  ODL ;
wire  ODM ;
wire  ODN ;
wire  ODO ;
wire  ODP ;
wire  OEA ;
wire  OEB ;
wire  OEC ;
wire  OED ;
wire  OEE ;
wire  OEF ;
wire  OEG ;
wire  OEH ;
wire  OEI ;
wire  OEJ ;
wire  OEK ;
wire  OEL ;
wire  OEM ;
wire  OEN ;
wire  OEO ;
wire  OEP ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OFE ;
wire  OFF ;
wire  OFG ;
wire  OFH ;
wire  OFI ;
wire  OFJ ;
wire  OFK ;
wire  OFL ;
wire  OFM ;
wire  OFN ;
wire  OFO ;
wire  OFP ;
wire  oga ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  okg ;
wire  okh ;
wire  oki ;
wire  okj ;
wire  okk ;
wire  okl ;
wire  okm ;
wire  okn ;
wire  oko ;
wire  okp ;
wire  OKQ ;
wire  okr ;
wire  oks ;
wire  okt ;
wire  ola ;
wire  OLB ;
wire  OLC ;
wire  OLD ;
wire  OLE ;
wire  olf ;
wire  olg ;
wire  OLH ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pai ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pan ;
wire  pao ;
wire  pap ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pco ;
wire  pcp ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pdj ;
wire  pdk ;
wire  pdl ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  pdp ;
wire  QAA ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  QAK ;
wire  QAL ;
wire  qam ;
wire  qan ;
wire  qao ;
wire  qap ;
wire  QAQ ;
wire  qat ;
wire  qba ;
wire  qbb ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qce ;
wire  qcf ;
wire  qcg ;
wire  qch ;
wire  qci ;
wire  qcj ;
wire  qck ;
wire  qcl ;
wire  qcm ;
wire  qcn ;
wire  qco ;
wire  qcp ;
wire  qcq ;
wire  qcr ;
wire  qcs ;
wire  qct ;
wire  qcu ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qdf ;
wire  qdg ;
wire  qdh ;
wire  qdi ;
wire  qdj ;
wire  qdk ;
wire  qdl ;
wire  qdm ;
wire  qdn ;
wire  qdo ;
wire  qea ;
wire  qeb ;
wire  qfa ;
wire  qfb ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  qge ;
wire  qgf ;
wire  qha ;
wire  qhb ;
wire  qhc ;
wire  qhd ;
wire  qhe ;
wire  qia ;
wire  qib ;
wire  qja ;
wire  qjb ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qkd ;
wire  qke ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  qma ;
wire  qmb ;
wire  qmc ;
wire  qmd ;
wire  QME ;
wire  qmf ;
wire  qmg ;
wire  QMH ;
wire  qmi ;
wire  qmj ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  qnd ;
wire  QOA ;
wire  QOB ;
wire  QOC ;
wire  qod ;
wire  qpa ;
wire  qpb ;
wire  qpc ;
wire  qpd ;
wire  qpe ;
wire  qpf ;
wire  qpg ;
wire  qph ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qqd ;
wire  qqe ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  qrf ;
wire  qrg ;
wire  qrh ;
wire  qri ;
wire  qrj ;
wire  qrk ;
wire  qrl ;
wire  qrm ;
wire  qrn ;
wire  qro ;
wire  qrp ;
wire  qsa ;
wire  qsb ;
wire  qsc ;
wire  qsd ;
wire  qse ;
wire  qsf ;
wire  qsg ;
wire  qsh ;
wire  qsi ;
wire  qsj ;
wire  qsk ;
wire  qsl ;
wire  qsm ;
wire  qsn ;
wire  qso ;
wire  qsp ;
wire  qta ;
wire  qtb ;
wire  qtc ;
wire  qtd ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qud ;
wire  QUE ;
wire  QUF ;
wire  qug ;
wire  quh ;
wire  qva ;
wire  qvb ;
wire  qvc ;
wire  saa ;
wire  sab ;
wire  sac ;
wire  sad ;
wire  sae ;
wire  saf ;
wire  sag ;
wire  sah ;
wire  sai ;
wire  saj ;
wire  sak ;
wire  sal ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tae ;
wire  TAE ;
wire  taf ;
wire  TAF ;
wire  tag ;
wire  TAG ;
wire  tah ;
wire  TAH ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tbe ;
wire  TBE ;
wire  tbf ;
wire  TBF ;
wire  tbg ;
wire  TBG ;
wire  tbh ;
wire  TBH ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tcg ;
wire  TCG ;
wire  tch ;
wire  TCH ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tde ;
wire  TDE ;
wire  tdf ;
wire  TDF ;
wire  tdg ;
wire  TDG ;
wire  tdh ;
wire  TDH ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tfa ;
wire  TFA ;
wire  tfb ;
wire  TFB ;
wire  tfc ;
wire  TFC ;
wire  tfd ;
wire  TFD ;
wire  tha ;
wire  THA ;
wire  thb ;
wire  THB ;
wire  thc ;
wire  THC ;
wire  tia ;
wire  TIA ;
wire  tib ;
wire  TIB ;
wire  tic ;
wire  TIC ;
wire  tid ;
wire  TID ;
wire  tie ;
wire  TIE ;
wire  tif ;
wire  TIF ;
wire  tig ;
wire  TIG ;
wire  tja ;
wire  TJA ;
wire  tjb ;
wire  TJB ;
wire  tjc ;
wire  TJC ;
wire  tjd ;
wire  TJD ;
wire  tje ;
wire  TJE ;
wire  tjf ;
wire  TJF ;
wire  tjg ;
wire  TJG ;
wire  tjh ;
wire  TJH ;
wire  tji ;
wire  TJI ;
wire  tjj ;
wire  TJJ ;
wire  tjk ;
wire  TJK ;
wire  tjl ;
wire  TJL ;
wire  tka ;
wire  TKA ;
wire  tkb ;
wire  TKB ;
wire  tkc ;
wire  TKC ;
wire  tkd ;
wire  TKD ;
wire  tla ;
wire  TLA ;
wire  tlb ;
wire  TLB ;
wire  tlc ;
wire  TLC ;
wire  tld ;
wire  TLD ;
wire  tma ;
wire  TMA ;
wire  tmb ;
wire  TMB ;
wire  tmc ;
wire  TMC ;
wire  tmd ;
wire  TMD ;
wire  tna ;
wire  TNA ;
wire  tnb ;
wire  TNB ;
wire  toa ;
wire  TOA ;
wire  tpa ;
wire  TPA ;
wire  tpb ;
wire  TPB ;
wire  tpc ;
wire  TPC ;
wire  tpd ;
wire  TPD ;
wire  tpe ;
wire  TPE ;
wire  tpf ;
wire  TPF ;
wire  tpg ;
wire  TPG ;
wire  tph ;
wire  TPH ;
wire  tpi ;
wire  TPI ;
wire  tpj ;
wire  TPJ ;
wire  tqa ;
wire  TQA ;
wire  tqb ;
wire  TQB ;
wire  tqc ;
wire  TQC ;
wire  tqd ;
wire  TQD ;
wire  tsa ;
wire  TSA ;
wire  tsb ;
wire  TSB ;
wire  tsc ;
wire  TSC ;
wire  tta ;
wire  TTA ;
wire  UAA ;
wire  UAB ;
wire  UAC ;
wire  UAD ;
wire  UAE ;
wire  UAF ;
wire  UAG ;
wire  UAH ;
wire  UAI ;
wire  UAJ ;
wire  UAK ;
wire  UAL ;
wire  UAM ;
wire  UAN ;
wire  UAO ;
wire  UAP ;
wire  UBA ;
wire  UBB ;
wire  UBC ;
wire  UBD ;
wire  UBE ;
wire  UBF ;
wire  UBG ;
wire  UBH ;
wire  UBI ;
wire  UBJ ;
wire  UBK ;
wire  UBL ;
wire  UBM ;
wire  UBN ;
wire  UBO ;
wire  UBP ;
wire  UCA ;
wire  UCB ;
wire  UCC ;
wire  UCD ;
wire  UCE ;
wire  UCF ;
wire  UCG ;
wire  UCH ;
wire  UCI ;
wire  UCJ ;
wire  UCK ;
wire  UCL ;
wire  UCM ;
wire  UCN ;
wire  UCO ;
wire  UCP ;
wire  UDA ;
wire  UDB ;
wire  UDC ;
wire  UDD ;
wire  UDE ;
wire  UDF ;
wire  UDG ;
wire  UDH ;
wire  UDI ;
wire  UDJ ;
wire  UDK ;
wire  UDL ;
wire  UDM ;
wire  UDN ;
wire  UDO ;
wire  UDP ;
wire  VAA ;
wire  VAB ;
wire  vac ;
wire  vad ;
wire  VBA ;
wire  VBB ;
wire  vbc ;
wire  vbd ;
wire  VCA ;
wire  VCB ;
wire  vcc ;
wire  vcd ;
wire  VDA ;
wire  VDB ;
wire  vdc ;
wire  vdd ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wai ;
wire  waj ;
wire  wak ;
wire  wal ;
wire  wam ;
wire  wan ;
wire  wao ;
wire  wap ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wbi ;
wire  wbj ;
wire  wbk ;
wire  wbl ;
wire  wbm ;
wire  wbn ;
wire  wbo ;
wire  wbp ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wci ;
wire  wcj ;
wire  wck ;
wire  wcl ;
wire  wcm ;
wire  wcn ;
wire  wco ;
wire  wcp ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wdi ;
wire  wdj ;
wire  wdk ;
wire  wdl ;
wire  wdm ;
wire  wdn ;
wire  wdo ;
wire  wdp ;
wire  xaa ;
wire  xab ;
wire  xac ;
wire  xad ;
wire  xae ;
wire  xaf ;
wire  xag ;
wire  xah ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign VAA = ~vaa;  //complement 
assign paa = ~PAA;  //complement 
assign xaa = ~XAA;  //complement 
assign VBA = ~vba;  //complement 
assign pai = ~PAI;  //complement 
assign FAA = QTA & BAA ; 
assign faa = ~FAA ; //complement 
assign FAI = QTA & BAI ; 
assign fai = ~FAI ;  //complement 
assign FBA = QTB & BBA ; 
assign fba = ~FBA ;  //complement 
assign FBI = QTB & BBI; 
assign fbi = ~FBI; 
assign VCA = ~vca;  //complement 
assign pba = ~PBA;  //complement 
assign BAA = ~baa;  //complement 
assign BAI = ~bai;  //complement 
assign VDA = ~vda;  //complement 
assign pbi = ~PBI;  //complement 
assign BBA = ~bba;  //complement 
assign BBI = ~bbi;  //complement 
assign vac = ~VAC;  //complement 
assign pca = ~PCA;  //complement 
assign BCA = ~bca;  //complement 
assign BCI = ~bci;  //complement 
assign vbc = ~VBC;  //complement 
assign pci = ~PCI;  //complement 
assign BDA = ~bda;  //complement 
assign BDI = ~bdi;  //complement 
assign vcc = ~VCC;  //complement 
assign pda = ~PDA;  //complement 
assign FCA = QTC & BCA ; 
assign fca = ~FCA ; //complement 
assign FCI = QTC & BCI ; 
assign fci = ~FCI ;  //complement 
assign vdc = ~VDC;  //complement 
assign pdi = ~PDI;  //complement 
assign FDA = QTD & BDA ; 
assign fda = ~FDA ; //complement 
assign FDI = QTD & BDI ; 
assign fdi = ~FDI ;  //complement 
assign JHA =  QVA  ; 
assign jha = ~JHA;  //complement  
assign lba = ~LBA;  //complement 
assign lbi = ~LBI;  //complement 
assign waa = ~WAA;  //complement 
assign wai = ~WAI;  //complement 
assign taa = qpa; 
assign TAA = ~taa; //complement 
assign tac = qpa; 
assign TAC = ~tac;  //complement 
assign tad = qpa; 
assign TAD = ~tad;  //complement 
assign tab = qpa; 
assign TAB = ~tab;  //complement 
assign wba = ~WBA;  //complement 
assign wbi = ~WBI;  //complement 
assign JQA =  QAJ & gaa & qrg  |  qaj & GAA & qrg  |  qaj & gaa & QRG  |  QAJ & GAA & QRG  ; 
assign jqa = ~JQA; //complement 
assign jqb =  QAJ & gaa & qrg  |  qaj & GAA & qrg  |  qaj & gaa & QRG  |  qaj & gaa & qrg  ; 
assign JQB = ~jqb;  //complement 
assign HAA = ~haa;  //complement 
assign HBA = ~hba;  //complement 
assign HCA = ~hca;  //complement 
assign HDA = ~hda;  //complement 
assign QAQ = ~qaq;  //complement 
assign qqe = ~QQE;  //complement 
assign qtd = ~QTD;  //complement 
assign qaj = ~QAJ;  //complement 
assign qrg = ~QRG;  //complement 
assign gaa = ~GAA;  //complement 
assign gai = ~GAI;  //complement 
assign HAI = ~hai;  //complement 
assign HBI = ~hbi;  //complement 
assign HCI = ~hci;  //complement 
assign HDI = ~hdi;  //complement 
assign qdd = ~QDD;  //complement 
assign TFA = QQE; 
assign tfa = ~TFA; //complement 
assign TFB = QQE; 
assign tfb = ~TFB;  //complement 
assign TFC = QQE; 
assign tfc = ~TFC;  //complement 
assign TFD = QQE; 
assign tfd = ~TFD;  //complement 
assign gba = ~GBA;  //complement 
assign gbi = ~GBI;  //complement 
assign taf = qpe; 
assign TAF = ~taf; //complement 
assign tag = qpe; 
assign TAG = ~tag;  //complement 
assign tah = qpe; 
assign TAH = ~tah;  //complement 
assign tae = qpe; 
assign TAE = ~tae;  //complement 
assign wca = ~WCA;  //complement 
assign wci = ~WCI;  //complement 
assign kaa = ~KAA;  //complement 
assign kai = ~KAI;  //complement 
assign qpa = ~QPA;  //complement 
assign qpe = ~QPE;  //complement 
assign wda = ~WDA;  //complement 
assign wdi = ~WDI;  //complement 
assign qre = ~QRE;  //complement 
assign qrf = ~QRF;  //complement 
assign qrh = ~QRH;  //complement 
assign qri = ~QRI;  //complement 
assign qrj = ~QRJ;  //complement 
assign qrk = ~QRK;  //complement 
assign qrl = ~QRL;  //complement 
assign qrm = ~QRM;  //complement 
assign JEA =  QME  ; 
assign jea = ~JEA;  //complement  
assign JFA =  LAA & QMI  ; 
assign jfa = ~JFA;  //complement 
assign OAA = ~oaa;  //complement 
assign OAI = ~oai;  //complement 
assign OEA = ~oea;  //complement 
assign gca = ~GCA;  //complement 
assign gci = ~GCI;  //complement 
assign eaa = ~EAA;  //complement 
assign eai = ~EAI;  //complement 
assign oga = ~OGA;  //complement 
assign naa = ~NAA;  //complement 
assign nai = ~NAI;  //complement 
assign lai = ~LAI;  //complement 
assign saa = ~SAA;  //complement 
assign sai = ~SAI;  //complement 
assign OBA = ~oba;  //complement 
assign OBI = ~obi;  //complement 
assign OEI = ~oei;  //complement 
assign nba = ~NBA;  //complement 
assign nbi = ~NBI;  //complement 
assign QAK = ~qak;  //complement 
assign QAL = ~qal;  //complement 
assign AAA = ~aaa;  //complement 
assign ABA = ~aba;  //complement 
assign ABI = ~abi;  //complement 
assign oka = ~OKA;  //complement 
assign nca = ~NCA;  //complement 
assign nci = ~NCI;  //complement 
assign tna =  qag  ; 
assign TNA = ~tna;  //complement 
assign tnb =  qag  ; 
assign TNB = ~tnb;  //complement 
assign AAI = ~aai;  //complement 
assign QAA = ~qaa;  //complement 
assign oki = ~OKI;  //complement 
assign nda = ~NDA;  //complement 
assign ndi = ~NDI;  //complement 
assign qan = ~QAN;  //complement 
assign qag = ~QAG;  //complement 
assign OCA = ~oca;  //complement 
assign OCI = ~oci;  //complement 
assign OFA = ~ofa;  //complement 
assign OKQ = ~okq;  //complement 
assign qap = ~QAP;  //complement 
assign gda = ~GDA;  //complement 
assign gdi = ~GDI;  //complement 
assign eba = ~EBA;  //complement 
assign ebi = ~EBI;  //complement 
assign oks = ~OKS;  //complement 
assign qac = ~QAC;  //complement 
assign qrn = ~QRN;  //complement 
assign qro = ~QRO;  //complement 
assign qrp = ~QRP;  //complement 
assign qsa = ~QSA;  //complement 
assign laa = ~LAA;  //complement 
assign jla =  qqd & qdd  ; 
assign JLA = ~jla;  //complement 
assign ODA = ~oda;  //complement 
assign ODI = ~odi;  //complement 
assign OFI = ~ofi;  //complement 
assign pab = ~PAB;  //complement 
assign xab = ~XAB;  //complement 
assign qma = ~QMA;  //complement 
assign paj = ~PAJ;  //complement 
assign FAB = QTA & BAB ; 
assign fab = ~FAB ; //complement 
assign FAJ = QTA & BAJ ; 
assign faj = ~FAJ ;  //complement 
assign FBB = QTB & BBB ; 
assign fbb = ~FBB ;  //complement 
assign FBJ = QTB & BBJ; 
assign fbj = ~FBJ; 
assign JAA =  QMA  ; 
assign jaa = ~JAA;  //complement  
assign JAB =  QMA & DAA  ; 
assign jab = ~JAB;  //complement 
assign pbb = ~PBB;  //complement 
assign BAB = ~bab;  //complement 
assign BAJ = ~baj;  //complement 
assign JAC =  QMA & DAA & DAB  ; 
assign jac = ~JAC;  //complement  
assign JAD =  QMA & DAA & DAB & DAC  ; 
assign jad = ~JAD;  //complement 
assign pbj = ~PBJ;  //complement 
assign BBB = ~bbb;  //complement 
assign BBJ = ~bbj;  //complement 
assign daa = ~DAA;  //complement 
assign pcb = ~PCB;  //complement 
assign BCB = ~bcb;  //complement 
assign BCJ = ~bcj;  //complement 
assign dab = ~DAB;  //complement 
assign pcj = ~PCJ;  //complement 
assign BDB = ~bdb;  //complement 
assign BDJ = ~bdj;  //complement 
assign dac = ~DAC;  //complement 
assign pdb = ~PDB;  //complement 
assign FCJ = QTC & BCJ ; 
assign fcj = ~FCJ ; //complement 
assign FCB = QTC & BCB ; 
assign fcb = ~FCB ;  //complement 
assign FDB = QTD & BDB ; 
assign fdb = ~FDB ;  //complement 
assign FDJ = QTD & BDJ; 
assign fdj = ~FDJ; 
assign dad = ~DAD;  //complement 
assign pdj = ~PDJ;  //complement 
assign JHB =  QVA & xaa  ; 
assign jhb = ~JHB;  //complement  
assign lbb = ~LBB;  //complement 
assign lbj = ~LBJ;  //complement 
assign wab = ~WAB;  //complement 
assign waj = ~WAJ;  //complement 
assign tba = qpb; 
assign TBA = ~tba; //complement 
assign tbb = qpb; 
assign TBB = ~tbb;  //complement 
assign tbc = qpb; 
assign TBC = ~tbc;  //complement 
assign tbd = qpb; 
assign TBD = ~tbd;  //complement 
assign wbb = ~WBB;  //complement 
assign wbj = ~WBJ;  //complement 
assign HAB = ~hab;  //complement 
assign HBB = ~hbb;  //complement 
assign HCB = ~hcb;  //complement 
assign HDB = ~hdb;  //complement 
assign gab = ~GAB;  //complement 
assign gaj = ~GAJ;  //complement 
assign HAJ = ~haj;  //complement 
assign HBJ = ~hbj;  //complement 
assign HCJ = ~hcj;  //complement 
assign HDJ = ~hdj;  //complement 
assign qce = ~QCE;  //complement 
assign gbb = ~GBB;  //complement 
assign gbj = ~GBJ;  //complement 
assign tbe = qpf; 
assign TBE = ~tbe; //complement 
assign tbf = qpf; 
assign TBF = ~tbf;  //complement 
assign tbg = qpf; 
assign TBG = ~tbg;  //complement 
assign tbh = qpf; 
assign TBH = ~tbh;  //complement 
assign wcb = ~WCB;  //complement 
assign wcj = ~WCJ;  //complement 
assign kab = ~KAB;  //complement 
assign kaj = ~KAJ;  //complement 
assign qpb = ~QPB;  //complement 
assign qpf = ~QPF;  //complement 
assign wdb = ~WDB;  //complement 
assign wdj = ~WDJ;  //complement 
assign TJG =  QIB  ; 
assign tjg = ~TJG;  //complement 
assign TJH =  QIA  ; 
assign tjh = ~TJH;  //complement 
assign qsb = ~QSB;  //complement 
assign qsc = ~QSC;  //complement 
assign qsd = ~QSD;  //complement 
assign qse = ~QSE;  //complement 
assign qsf = ~QSF;  //complement 
assign qsg = ~QSG;  //complement 
assign qsh = ~QSH;  //complement 
assign qsi = ~QSI;  //complement 
assign JEB =  QME & lba  ; 
assign jeb = ~JEB;  //complement  
assign JFB =  LAB & QMI  ; 
assign jfb = ~JFB;  //complement 
assign OAB = ~oab;  //complement 
assign OAJ = ~oaj;  //complement 
assign OEB = ~oeb;  //complement 
assign tie =  qca & qda & qua  ; 
assign TIE = ~tie;  //complement 
assign tsb =  qba  ; 
assign TSB = ~tsb;  //complement 
assign gcb = ~GCB;  //complement 
assign gcj = ~GCJ;  //complement 
assign eab = ~EAB;  //complement 
assign eaj = ~EAJ;  //complement 
assign OGB = ~ogb;  //complement 
assign nab = ~NAB;  //complement 
assign naj = ~NAJ;  //complement 
assign sab = ~SAB;  //complement 
assign saj = ~SAJ;  //complement 
assign OBB = ~obb;  //complement 
assign OBJ = ~obj;  //complement 
assign OEJ = ~oej;  //complement 
assign OLB = ~olb;  //complement 
assign nbb = ~NBB;  //complement 
assign nbj = ~NBJ;  //complement 
assign TOA =  QBB  ; 
assign toa = ~TOA;  //complement 
assign TSA =  qak & qal & qba  ; 
assign tsa = ~TSA;  //complement 
assign tsc =  qak & qal & qba  ; 
assign TSC = ~tsc;  //complement 
assign AAB = ~aab;  //complement 
assign ABB = ~abb;  //complement 
assign ABJ = ~abj;  //complement 
assign okb = ~OKB;  //complement 
assign ncb = ~NCB;  //complement 
assign ncj = ~NCJ;  //complement 
assign JKB =  cam & cal & cak & CAJ  ; 
assign jkb = ~JKB;  //complement  
assign JKI =  CAM & cbl & cbk & cbj  ; 
assign jki = ~JKI;  //complement 
assign AAJ = ~aaj;  //complement 
assign CAJ = ~caj;  //complement 
assign CBJ = ~cbj;  //complement 
assign okj = ~OKJ;  //complement 
assign ndb = ~NDB;  //complement 
assign ndj = ~NDJ;  //complement 
assign qia = ~QIA;  //complement 
assign qba = ~QBA;  //complement 
assign OCB = ~ocb;  //complement 
assign OCJ = ~ocj;  //complement 
assign OFB = ~ofb;  //complement 
assign OLD = ~old;  //complement 
assign qbb = ~QBB;  //complement 
assign qib = ~QIB;  //complement 
assign gdb = ~GDB;  //complement 
assign gdj = ~GDJ;  //complement 
assign ebb = ~EBB;  //complement 
assign ebj = ~EBJ;  //complement 
assign qsj = ~QSJ;  //complement 
assign qsk = ~QSK;  //complement 
assign qsl = ~QSL;  //complement 
assign qsm = ~QSM;  //complement 
assign lab = ~LAB;  //complement 
assign laj = ~LAJ;  //complement 
assign ODB = ~odb;  //complement 
assign ODJ = ~odj;  //complement 
assign OFJ = ~ofj;  //complement 
assign pac = ~PAC;  //complement 
assign xac = ~XAC;  //complement 
assign qmb = ~QMB;  //complement 
assign pak = ~PAK;  //complement 
assign FAC = QTA & BAC ; 
assign fac = ~FAC ; //complement 
assign FAK = QTA & BAK ; 
assign fak = ~FAK ;  //complement 
assign FBC = QTB & BBC ; 
assign fbc = ~FBC ;  //complement 
assign FBK = QTB & BBK; 
assign fbk = ~FBK; 
assign JBA =  QMB  ; 
assign jba = ~JBA;  //complement  
assign JBB =  QMB & DBA  ; 
assign jbb = ~JBB;  //complement 
assign pbc = ~PBC;  //complement 
assign BAC = ~bac;  //complement 
assign BAK = ~bak;  //complement 
assign JBC =  QMB & DBA & DBB  ; 
assign jbc = ~JBC;  //complement  
assign JBD =  QMB & DBA & DBB & DBC  ; 
assign jbd = ~JBD;  //complement 
assign pbk = ~PBK;  //complement 
assign BBC = ~bbc;  //complement 
assign BBK = ~bbk;  //complement 
assign dba = ~DBA;  //complement 
assign pcc = ~PCC;  //complement 
assign BCC = ~bcc;  //complement 
assign BCK = ~bck;  //complement 
assign dbb = ~DBB;  //complement 
assign pck = ~PCK;  //complement 
assign BDC = ~bdc;  //complement 
assign BDK = ~bdk;  //complement 
assign dbc = ~DBC;  //complement 
assign pdc = ~PDC;  //complement 
assign FDD = QTD & BDD ; 
assign fdd = ~FDD ; //complement 
assign FDC = QTD & BDC ; 
assign fdc = ~FDC ;  //complement 
assign FDK = QTD & BDK ; 
assign fdk = ~FDK ;  //complement 
assign FDL = QTD & BDL; 
assign fdl = ~FDL; 
assign FCG = QTC & BCH ; 
assign fcg = ~FCG ; //complement 
assign FCK = QTC & BCK ; 
assign fck = ~FCK ;  //complement 
assign FCC = QTC & BCC ; 
assign fcc = ~FCC ;  //complement 
assign dbd = ~DBD;  //complement 
assign pdk = ~PDK;  //complement 
assign JHC =  QVA & xaa & xab  ; 
assign jhc = ~JHC;  //complement  
assign qnd = ~QND;  //complement 
assign lbc = ~LBC;  //complement 
assign lbk = ~LBK;  //complement 
assign qcg = ~QCG;  //complement 
assign qch = ~QCH;  //complement 
assign qci = ~QCI;  //complement 
assign wac = ~WAC;  //complement 
assign wak = ~WAK;  //complement 
assign qct = ~QCT;  //complement 
assign qcu = ~QCU;  //complement 
assign tca = qpc; 
assign TCA = ~tca; //complement 
assign tcb = qpc; 
assign TCB = ~tcb;  //complement 
assign tcc = qpc; 
assign TCC = ~tcc;  //complement 
assign tcd = qpc; 
assign TCD = ~tcd;  //complement 
assign wbc = ~WBC;  //complement 
assign wbk = ~WBK;  //complement 
assign qcn = ~QCN;  //complement 
assign qcq = ~QCQ;  //complement 
assign qcr = ~QCR;  //complement 
assign qcs = ~QCS;  //complement 
assign HAC = ~hac;  //complement 
assign HBC = ~hbc;  //complement 
assign HCC = ~hcc;  //complement 
assign HDC = ~hdc;  //complement 
assign qcb = ~QCB;  //complement 
assign qcf = ~QCF;  //complement 
assign qcc = ~QCC;  //complement 
assign qcj = ~QCJ;  //complement 
assign qcl = ~QCL;  //complement 
assign qcm = ~QCM;  //complement 
assign gac = ~GAC;  //complement 
assign gak = ~GAK;  //complement 
assign HAK = ~hak;  //complement 
assign HBK = ~hbk;  //complement 
assign HCK = ~hck;  //complement 
assign HDK = ~hdk;  //complement 
assign qco = ~QCO;  //complement 
assign qck = ~QCK;  //complement 
assign qcp = ~QCP;  //complement 
assign gbc = ~GBC;  //complement 
assign gbk = ~GBK;  //complement 
assign tce = qpg; 
assign TCE = ~tce; //complement 
assign tcf = qpg; 
assign TCF = ~tcf;  //complement 
assign tcg = qpg; 
assign TCG = ~tcg;  //complement 
assign tch = qpg; 
assign TCH = ~tch;  //complement 
assign wcc = ~WCC;  //complement 
assign wck = ~WCK;  //complement 
assign kac = ~KAC;  //complement 
assign kak = ~KAK;  //complement 
assign qpc = ~QPC;  //complement 
assign qpg = ~QPG;  //complement 
assign wdc = ~WDC;  //complement 
assign wdk = ~WDK;  //complement 
assign jlb =  qcc & qcf & qcr  ; 
assign JLB = ~jlb;  //complement 
assign TJE =  QJB  ; 
assign tje = ~TJE;  //complement 
assign TJF =  QJA  ; 
assign tjf = ~TJF;  //complement 
assign qkc = ~QKC;  //complement 
assign JEC =  QME & lba & lbb  ; 
assign jec = ~JEC;  //complement  
assign JFC =  LAC & QMI  ; 
assign jfc = ~JFC;  //complement 
assign OAC = ~oac;  //complement 
assign OAK = ~oak;  //complement 
assign OEC = ~oec;  //complement 
assign TPD = QOC; 
assign tpd = ~TPD; //complement 
assign TPC = QOC; 
assign tpc = ~TPC;  //complement 
assign TPE = QAI; 
assign tpe = ~TPE;  //complement 
assign TPF = QAI; 
assign tpf = ~TPF;  //complement 
assign gcc = ~GCC;  //complement 
assign gck = ~GCK;  //complement 
assign eac = ~EAC;  //complement 
assign eak = ~EAK;  //complement 
assign OGC = ~ogc;  //complement 
assign nac = ~NAC;  //complement 
assign nak = ~NAK;  //complement 
assign lac = ~LAC;  //complement 
assign sac = ~SAC;  //complement 
assign OBC = ~obc;  //complement 
assign OBK = ~obk;  //complement 
assign OEK = ~oek;  //complement 
assign qjb = ~QJB;  //complement 
assign nbc = ~NBC;  //complement 
assign nbk = ~NBK;  //complement 
assign AAC = ~aac;  //complement 
assign ABC = ~abc;  //complement 
assign ABK = ~abk;  //complement 
assign okc = ~OKC;  //complement 
assign ncc = ~NCC;  //complement 
assign nck = ~NCK;  //complement 
assign JKC =  cam & cal & CAK & caj  ; 
assign jkc = ~JKC;  //complement  
assign JKJ =  CAM & cbl & cbk & CBJ  ; 
assign jkj = ~JKJ;  //complement 
assign AAK = ~aak;  //complement 
assign CAK = ~cak;  //complement 
assign CBK = ~cbk;  //complement 
assign okk = ~OKK;  //complement 
assign ndc = ~NDC;  //complement 
assign ndk = ~NDK;  //complement 
assign qca = ~QCA;  //complement 
assign qja = ~QJA;  //complement 
assign sak = ~SAK;  //complement 
assign OCC = ~occ;  //complement 
assign OCK = ~ock;  //complement 
assign OFC = ~ofc;  //complement 
assign OLC = ~olc;  //complement 
assign gdc = ~GDC;  //complement 
assign gdk = ~GDK;  //complement 
assign ebc = ~EBC;  //complement 
assign ebk = ~EBK;  //complement 
assign ODC = ~odc;  //complement 
assign ODK = ~odk;  //complement 
assign OFK = ~ofk;  //complement 
assign UAA = ~uaa;  //complement 
assign UAB = ~uab;  //complement 
assign UAC = ~uac;  //complement 
assign UAD = ~uad;  //complement 
assign pad = ~PAD;  //complement 
assign xad = ~XAD;  //complement 
assign UAI = ~uai;  //complement 
assign UAJ = ~uaj;  //complement 
assign UAK = ~uak;  //complement 
assign UAL = ~ual;  //complement 
assign pal = ~PAL;  //complement 
assign FBD = QTB & BBD ; 
assign fbd = ~FBD ; //complement 
assign FBL = QTB & BBL ; 
assign fbl = ~FBL ;  //complement 
assign FAD = QTA & BAD ; 
assign fad = ~FAD ;  //complement 
assign FAL = QTA & BAL; 
assign fal = ~FAL; 
assign UBA = ~uba;  //complement 
assign UBB = ~ubb;  //complement 
assign UBC = ~ubc;  //complement 
assign UBD = ~ubd;  //complement 
assign pbd = ~PBD;  //complement 
assign BAD = ~bad;  //complement 
assign BAL = ~bal;  //complement 
assign UBI = ~ubi;  //complement 
assign UBJ = ~ubj;  //complement 
assign UBK = ~ubk;  //complement 
assign UBL = ~ubl;  //complement 
assign pbl = ~PBL;  //complement 
assign BBD = ~bbd;  //complement 
assign BBL = ~bbl;  //complement 
assign UCA = ~uca;  //complement 
assign UCB = ~ucb;  //complement 
assign UCC = ~ucc;  //complement 
assign UCD = ~ucd;  //complement 
assign pcd = ~PCD;  //complement 
assign BCD = ~bcd;  //complement 
assign BCL = ~bcl;  //complement 
assign UCI = ~uci;  //complement 
assign UCJ = ~ucj;  //complement 
assign UCK = ~uck;  //complement 
assign UCL = ~ucl;  //complement 
assign pcl = ~PCL;  //complement 
assign BDD = ~bdd;  //complement 
assign BDL = ~bdl;  //complement 
assign UDA = ~uda;  //complement 
assign UDB = ~udb;  //complement 
assign UDC = ~udc;  //complement 
assign UDD = ~udd;  //complement 
assign pdd = ~PDD;  //complement 
assign FCD = QTC & BCD ; 
assign fcd = ~FCD ; //complement 
assign FCL = QTC & BCL ; 
assign fcl = ~FCL ;  //complement 
assign UDI = ~udi;  //complement 
assign UDJ = ~udj;  //complement 
assign UDK = ~udk;  //complement 
assign UDL = ~udl;  //complement 
assign pdl = ~PDL;  //complement 
assign JHD =  QVA & xaa & xab & xac  ; 
assign jhd = ~JHD;  //complement  
assign JIA =  xaa & xab & xac & xad  ; 
assign jia = ~JIA;  //complement 
assign lbd = ~LBD;  //complement 
assign lbl = ~LBL;  //complement 
assign JOA =  QHD  ; 
assign joa = ~JOA;  //complement 
assign wad = ~WAD;  //complement 
assign wal = ~WAL;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign qdf = ~QDF;  //complement 
assign qdg = ~QDG;  //complement 
assign tda = qpd; 
assign TDA = ~tda; //complement 
assign tdb = qpd; 
assign TDB = ~tdb;  //complement 
assign tdc = qpd; 
assign TDC = ~tdc;  //complement 
assign tdd = qpd; 
assign TDD = ~tdd;  //complement 
assign wbd = ~WBD;  //complement 
assign wbl = ~WBL;  //complement 
assign qdh = ~QDH;  //complement 
assign qdl = ~QDL;  //complement 
assign qdm = ~QDM;  //complement 
assign qdn = ~QDN;  //complement 
assign HAD = ~had;  //complement 
assign HBD = ~hbd;  //complement 
assign HCD = ~hcd;  //complement 
assign HDD = ~hdd;  //complement 
assign qdo = ~QDO;  //complement 
assign qde = ~QDE;  //complement 
assign gad = ~GAD;  //complement 
assign gal = ~GAL;  //complement 
assign HAL = ~hal;  //complement 
assign HBL = ~hbl;  //complement 
assign HCL = ~hcl;  //complement 
assign HDL = ~hdl;  //complement 
assign qdj = ~QDJ;  //complement 
assign qdk = ~QDK;  //complement 
assign qmg = ~QMG;  //complement 
assign gbd = ~GBD;  //complement 
assign gbl = ~GBL;  //complement 
assign tde = qph; 
assign TDE = ~tde; //complement 
assign tdf = qph; 
assign TDF = ~tdf;  //complement 
assign tdg = qph; 
assign TDG = ~tdg;  //complement 
assign tdh = qph; 
assign TDH = ~tdh;  //complement 
assign qdi = ~QDI;  //complement 
assign wcd = ~WCD;  //complement 
assign wcl = ~WCL;  //complement 
assign kad = ~KAD;  //complement 
assign kal = ~KAL;  //complement 
assign qpd = ~QPD;  //complement 
assign qph = ~QPH;  //complement 
assign wdd = ~WDD;  //complement 
assign wdl = ~WDL;  //complement 
assign jlc =  qdc & qdi & qdo  ; 
assign JLC = ~jlc;  //complement 
assign qra = ~QRA;  //complement 
assign qrb = ~QRB;  //complement 
assign qrc = ~QRC;  //complement 
assign qrd = ~QRD;  //complement 
assign qsn = ~QSN;  //complement 
assign qso = ~QSO;  //complement 
assign qsp = ~QSP;  //complement 
assign JED =  QME & lba & lbb & lbc  ; 
assign jed = ~JED;  //complement  
assign JFD =  LAD & QMI  ; 
assign jfd = ~JFD;  //complement 
assign OGE = ~oge;  //complement 
assign OAD = ~oad;  //complement 
assign OAL = ~oal;  //complement 
assign OED = ~oed;  //complement 
assign tpg = qah; 
assign TPG = ~tpg; //complement 
assign tph = qah; 
assign TPH = ~tph;  //complement 
assign tpi = qah; 
assign TPI = ~tpi;  //complement 
assign tpj = qah; 
assign TPJ = ~tpj;  //complement 
assign gcd = ~GCD;  //complement 
assign gcl = ~GCL;  //complement 
assign ead = ~EAD;  //complement 
assign eal = ~EAL;  //complement 
assign OGD = ~ogd;  //complement 
assign ohb = ~OHB;  //complement 
assign nad = ~NAD;  //complement 
assign nal = ~NAL;  //complement 
assign lad = ~LAD;  //complement 
assign sad = ~SAD;  //complement 
assign OBD = ~obd;  //complement 
assign OBL = ~obl;  //complement 
assign OEL = ~oel;  //complement 
assign nbd = ~NBD;  //complement 
assign nbl = ~NBL;  //complement 
assign oha = ~OHA;  //complement 
assign qah = ~QAH;  //complement 
assign AAD = ~aad;  //complement 
assign ABD = ~abd;  //complement 
assign ABL = ~abl;  //complement 
assign OLE = ~ole;  //complement 
assign okd = ~OKD;  //complement 
assign ncd = ~NCD;  //complement 
assign ncl = ~NCL;  //complement 
assign JKD =  cam & cal & CAK & CAJ  ; 
assign jkd = ~JKD;  //complement  
assign JKK =  CAM & cbl & CBK & cbj  ; 
assign jkk = ~JKK;  //complement 
assign AAL = ~aal;  //complement 
assign CAL = ~cal;  //complement 
assign CBL = ~cbl;  //complement 
assign okl = ~OKL;  //complement 
assign ndd = ~NDD;  //complement 
assign ndl = ~NDL;  //complement 
assign qda = ~QDA;  //complement 
assign qka = ~QKA;  //complement 
assign sal = ~SAL;  //complement 
assign OCD = ~ocd;  //complement 
assign OCL = ~ocl;  //complement 
assign OFD = ~ofd;  //complement 
assign qaf = ~QAF;  //complement 
assign TPA = qod & qai ; 
assign tpa = ~TPA ; //complement 
assign TPB = qod & qai ; 
assign tpb = ~TPB ;  //complement 
assign gdd = ~GDD;  //complement 
assign gdl = ~GDL;  //complement 
assign ebd = ~EBD;  //complement 
assign ebl = ~EBL;  //complement 
assign ola = ~OLA;  //complement 
assign qai = ~QAI;  //complement 
assign ODD = ~odd;  //complement 
assign ODL = ~odl;  //complement 
assign OFL = ~ofl;  //complement 
assign UAE = ~uae;  //complement 
assign UAF = ~uaf;  //complement 
assign UAG = ~uag;  //complement 
assign UAH = ~uah;  //complement 
assign pae = ~PAE;  //complement 
assign xae = ~XAE;  //complement 
assign UAM = ~uam;  //complement 
assign UAN = ~uan;  //complement 
assign UAO = ~uao;  //complement 
assign UAP = ~uap;  //complement 
assign pam = ~PAM;  //complement 
assign FAE = QTA & BAE ; 
assign fae = ~FAE ; //complement 
assign FAM = QTA & BAM ; 
assign fam = ~FAM ;  //complement 
assign FBE = QTB & BBE ; 
assign fbe = ~FBE ;  //complement 
assign FBM = QTB & BBM; 
assign fbm = ~FBM; 
assign UBE = ~ube;  //complement 
assign UBF = ~ubf;  //complement 
assign UBG = ~ubg;  //complement 
assign UBH = ~ubh;  //complement 
assign pbe = ~PBE;  //complement 
assign BAE = ~bae;  //complement 
assign BAM = ~bam;  //complement 
assign UBM = ~ubm;  //complement 
assign UBN = ~ubn;  //complement 
assign UBO = ~ubo;  //complement 
assign UBP = ~ubp;  //complement 
assign pbm = ~PBM;  //complement 
assign BBE = ~bbe;  //complement 
assign BBM = ~bbm;  //complement 
assign UCE = ~uce;  //complement 
assign UCF = ~ucf;  //complement 
assign UCG = ~ucg;  //complement 
assign UCH = ~uch;  //complement 
assign pce = ~PCE;  //complement 
assign BCE = ~bce;  //complement 
assign BCM = ~bcm;  //complement 
assign UCM = ~ucm;  //complement 
assign UCN = ~ucn;  //complement 
assign UCO = ~uco;  //complement 
assign UCP = ~ucp;  //complement 
assign pcm = ~PCM;  //complement 
assign BDE = ~bde;  //complement 
assign BDM = ~bdm;  //complement 
assign UDE = ~ude;  //complement 
assign UDF = ~udf;  //complement 
assign UDG = ~udg;  //complement 
assign UDH = ~udh;  //complement 
assign wde = ~WDE;  //complement 
assign FCE = QTC & BCE ; 
assign fce = ~FCE ; //complement 
assign FCM = QTC & BCM ; 
assign fcm = ~FCM ;  //complement 
assign FDM = QTD & BDM ; 
assign fdm = ~FDM ;  //complement 
assign FDE = QTD & BDE; 
assign fde = ~FDE; 
assign UDM = ~udm;  //complement 
assign UDN = ~udn;  //complement 
assign UDO = ~udo;  //complement 
assign UDP = ~udp;  //complement 
assign pdm = ~PDM;  //complement 
assign TIA = QQA; 
assign tia = ~TIA; //complement 
assign TIB = QQA; 
assign tib = ~TIB;  //complement 
assign TIC = QQA; 
assign tic = ~TIC;  //complement 
assign TID = QQA; 
assign tid = ~TID;  //complement 
assign JHE =  QVB  ; 
assign jhe = ~JHE;  //complement  
assign qna = ~QNA;  //complement 
assign lbe = ~LBE;  //complement 
assign lbm = ~LBM;  //complement 
assign wae = ~WAE;  //complement 
assign wam = ~WAM;  //complement 
assign job =  qcl & qdg  ; 
assign JOB = ~job;  //complement 
assign tja =  qcn  ; 
assign TJA = ~tja;  //complement 
assign tjb =  qcm  ; 
assign TJB = ~tjb;  //complement 
assign qqa = ~QQA;  //complement 
assign wbe = ~WBE;  //complement 
assign wbm = ~WBM;  //complement 
assign tjc =  qcl  ; 
assign TJC = ~tjc;  //complement 
assign tjd =  qck  ; 
assign TJD = ~tjd;  //complement 
assign HAE = ~hae;  //complement 
assign HBE = ~hbe;  //complement 
assign HCE = ~hce;  //complement 
assign HDE = ~hde;  //complement 
assign gae = ~GAE;  //complement 
assign gam = ~GAM;  //complement 
assign HAM = ~ham;  //complement 
assign HBM = ~hbm;  //complement 
assign HCM = ~hcm;  //complement 
assign HDM = ~hdm;  //complement 
assign qqd = ~QQD;  //complement 
assign qae = ~QAE;  //complement 
assign qqc = ~QQC;  //complement 
assign gbe = ~GBE;  //complement 
assign gbm = ~GBM;  //complement 
assign tif =  qqa  ; 
assign TIF = ~tif;  //complement 
assign tqa =  qao & qae  ; 
assign TQA = ~tqa;  //complement 
assign tqb =  qqa  ; 
assign TQB = ~tqb;  //complement 
assign wce = ~WCE;  //complement 
assign wcm = ~WCM;  //complement 
assign kae = ~KAE;  //complement 
assign kam = ~KAM;  //complement 
assign qmj = ~QMJ;  //complement 
assign qao = ~QAO;  //complement 
assign wdm = ~WDM;  //complement 
assign TJI =  QEB  ; 
assign tji = ~TJI;  //complement 
assign TJL =  QAM  ; 
assign tjl = ~TJL;  //complement 
assign pde = ~PDE;  //complement 
assign JEE =  QME & lba & lbb & lbc & lbd  ; 
assign jee = ~JEE;  //complement  
assign JFE =  LAE & QMI  ; 
assign jfe = ~JFE;  //complement 
assign OAE = ~oae;  //complement 
assign OAM = ~oam;  //complement 
assign OEE = ~oee;  //complement 
assign tig =  qcb & qdb & qub  ; 
assign TIG = ~tig;  //complement 
assign eae = ~EAE;  //complement 
assign eam = ~EAM;  //complement 
assign jna =  qcu & qgf & qhe & qbb & qea & qfa  ; 
assign JNA = ~jna;  //complement  
assign jnb =  qia & qja & qka & qla  ; 
assign JNB = ~jnb;  //complement 
assign nae = ~NAE;  //complement 
assign nam = ~NAM;  //complement 
assign lae = ~LAE;  //complement 
assign sae = ~SAE;  //complement 
assign OBE = ~obe;  //complement 
assign OBM = ~obm;  //complement 
assign OEM = ~oem;  //complement 
assign ohg = ~OHG;  //complement 
assign nbe = ~NBE;  //complement 
assign nbm = ~NBM;  //complement 
assign THA = qqd & qan ; 
assign tha = ~THA ; //complement 
assign THB = qqd & qan ; 
assign thb = ~THB ;  //complement 
assign AAE = ~aae;  //complement 
assign ABE = ~abe;  //complement 
assign ABM = ~abm;  //complement 
assign oke = ~OKE;  //complement 
assign nce = ~NCE;  //complement 
assign ncm = ~NCM;  //complement 
assign JKE =  cam & CAL & cak & caj  ; 
assign jke = ~JKE;  //complement  
assign JKL =  CAM & cbl & CBK & CBJ  ; 
assign jkl = ~JKL;  //complement 
assign AAM = ~aam;  //complement 
assign CAM = ~cam;  //complement 
assign CBM = ~cbm;  //complement 
assign okm = ~OKM;  //complement 
assign nde = ~NDE;  //complement 
assign ndm = ~NDM;  //complement 
assign qea = ~QEA;  //complement 
assign qla = ~QLA;  //complement 
assign OCE = ~oce;  //complement 
assign OCM = ~ocm;  //complement 
assign OFE = ~ofe;  //complement 
assign qeb = ~QEB;  //complement 
assign gde = ~GDE;  //complement 
assign gdm = ~GDM;  //complement 
assign ebe = ~EBE;  //complement 
assign ebm = ~EBM;  //complement 
assign ohd = ~OHD;  //complement 
assign ohe = ~OHE;  //complement 
assign ohf = ~OHF;  //complement 
assign gce = ~GCE;  //complement 
assign gcm = ~GCM;  //complement 
assign ODE = ~ode;  //complement 
assign ODM = ~odm;  //complement 
assign OFM = ~ofm;  //complement 
assign JCB =  QMC & DCA  ; 
assign jcb = ~JCB;  //complement  
assign paf = ~PAF;  //complement 
assign xaf = ~XAF;  //complement 
assign qmc = ~QMC;  //complement 
assign pan = ~PAN;  //complement 
assign FAF = QTA & BAF ; 
assign faf = ~FAF ; //complement 
assign FAN = QTA & BAN ; 
assign fan = ~FAN ;  //complement 
assign FBF = QTB & BBF ; 
assign fbf = ~FBF ;  //complement 
assign FBN = QTB & BBN; 
assign fbn = ~FBN; 
assign JCA =  QMC  ; 
assign jca = ~JCA;  //complement  
assign pbf = ~PBF;  //complement 
assign BAF = ~baf;  //complement 
assign BAN = ~ban;  //complement 
assign JCC =  QMC & DCA & DCB  ; 
assign jcc = ~JCC;  //complement  
assign JCD =  QMC & DCA & DCB & DCC  ; 
assign jcd = ~JCD;  //complement 
assign pbn = ~PBN;  //complement 
assign BBF = ~bbf;  //complement 
assign BBN = ~bbn;  //complement 
assign dca = ~DCA;  //complement 
assign pcf = ~PCF;  //complement 
assign BCF = ~bcf;  //complement 
assign BCN = ~bcn;  //complement 
assign dcb = ~DCB;  //complement 
assign pcn = ~PCN;  //complement 
assign BDF = ~bdf;  //complement 
assign BDN = ~bdn;  //complement 
assign dcc = ~DCC;  //complement 
assign pdf = ~PDF;  //complement 
assign FCF = QTC & BCF ; 
assign fcf = ~FCF ; //complement 
assign FCN = QTC & BCN ; 
assign fcn = ~FCN ;  //complement 
assign dcd = ~DCD;  //complement 
assign pdn = ~PDN;  //complement 
assign FDF = QTD & BDF ; 
assign fdf = ~FDF ; //complement 
assign FDN = QTD & BDN ; 
assign fdn = ~FDN ;  //complement 
assign JHF =  QVB & xae  ; 
assign jhf = ~JHF;  //complement  
assign qnb = ~QNB;  //complement 
assign lbf = ~LBF;  //complement 
assign lbn = ~LBN;  //complement 
assign qvb = ~QVB;  //complement 
assign qvc = ~QVC;  //complement 
assign waf = ~WAF;  //complement 
assign wan = ~WAN;  //complement 
assign qub = ~QUB;  //complement 
assign qva = ~QVA;  //complement 
assign wbf = ~WBF;  //complement 
assign wbn = ~WBN;  //complement 
assign HAF = ~haf;  //complement 
assign HBF = ~hbf;  //complement 
assign HCF = ~hcf;  //complement 
assign HDF = ~hdf;  //complement 
assign TTA =  QUB  ; 
assign tta = ~TTA;  //complement 
assign quc = ~QUC;  //complement 
assign qug = ~QUG;  //complement 
assign gaf = ~GAF;  //complement 
assign gan = ~GAN;  //complement 
assign HAN = ~han;  //complement 
assign HBN = ~hbn;  //complement 
assign HCN = ~hcn;  //complement 
assign HDN = ~hdn;  //complement 
assign qud = ~QUD;  //complement 
assign QUE = ~que;  //complement 
assign QUF = ~quf;  //complement 
assign gbf = ~GBF;  //complement 
assign gbn = ~GBN;  //complement 
assign jld =  qhc & quc  ; 
assign JLD = ~jld;  //complement 
assign tqc =  qao & qae & qhc  ; 
assign TQC = ~tqc;  //complement 
assign qam = ~QAM;  //complement 
assign wcf = ~WCF;  //complement 
assign wcn = ~WCN;  //complement 
assign kaf = ~KAF;  //complement 
assign kan = ~KAN;  //complement 
assign wdf = ~WDF;  //complement 
assign wdn = ~WDN;  //complement 
assign JEF =  QME & lba & lbb & lbc & lbd & lbe  ; 
assign jef = ~JEF;  //complement  
assign JFF =  LAF & QMI  ; 
assign jff = ~JFF;  //complement 
assign OAF = ~oaf;  //complement 
assign OAN = ~oan;  //complement 
assign OEF = ~oef;  //complement 
assign gcf = ~GCF;  //complement 
assign gcn = ~GCN;  //complement 
assign eaf = ~EAF;  //complement 
assign ean = ~EAN;  //complement 
assign OGF = ~ogf;  //complement 
assign naf = ~NAF;  //complement 
assign nan = ~NAN;  //complement 
assign laf = ~LAF;  //complement 
assign saf = ~SAF;  //complement 
assign OBF = ~obf;  //complement 
assign OBN = ~obn;  //complement 
assign OEN = ~oen;  //complement 
assign quh = ~QUH;  //complement 
assign nbf = ~NBF;  //complement 
assign nbn = ~NBN;  //complement 
assign ohc = ~OHC;  //complement 
assign AAF = ~aaf;  //complement 
assign ABF = ~abf;  //complement 
assign ABN = ~abn;  //complement 
assign okf = ~OKF;  //complement 
assign ncf = ~NCF;  //complement 
assign ncn = ~NCN;  //complement 
assign JKA =  cbm & cbl & cbk & cbj  ; 
assign jka = ~JKA;  //complement  
assign JKF =  cam & CAL & cak & CAJ  ; 
assign jkf = ~JKF;  //complement 
assign AAN = ~aan;  //complement 
assign CAN = ~can;  //complement 
assign okn = ~OKN;  //complement 
assign ndf = ~NDF;  //complement 
assign ndn = ~NDN;  //complement 
assign qfa = ~QFA;  //complement 
assign qfb = ~QFB;  //complement 
assign OCF = ~ocf;  //complement 
assign OCN = ~ocn;  //complement 
assign OFF = ~off;  //complement 
assign OLH = ~olh;  //complement 
assign TJJ =  QFB  ; 
assign tjj = ~TJJ;  //complement 
assign TJK =  QFA  ; 
assign tjk = ~TJK;  //complement 
assign gdf = ~GDF;  //complement 
assign gdn = ~GDN;  //complement 
assign ebf = ~EBF;  //complement 
assign ebn = ~EBN;  //complement 
assign ODF = ~odf;  //complement 
assign ODN = ~odn;  //complement 
assign OFN = ~ofn;  //complement 
assign pag = ~PAG;  //complement 
assign xag = ~XAG;  //complement 
assign qmd = ~QMD;  //complement 
assign pao = ~PAO;  //complement 
assign FAG = QTA & BAG ; 
assign fag = ~FAG ; //complement 
assign FAO = QTA & BAO ; 
assign fao = ~FAO ;  //complement 
assign FBG = QTB & BBG ; 
assign fbg = ~FBG ;  //complement 
assign FBO = QTB & BBO; 
assign fbo = ~FBO; 
assign JDA =  QMD  ; 
assign jda = ~JDA;  //complement  
assign JDB =  QMD & DDA  ; 
assign jdb = ~JDB;  //complement 
assign pbg = ~PBG;  //complement 
assign BAG = ~bag;  //complement 
assign BAO = ~bao;  //complement 
assign JDC =  QMD & DDA & DDB  ; 
assign jdc = ~JDC;  //complement  
assign JDD =  QMD & DDA & DDB & DDC  ; 
assign jdd = ~JDD;  //complement 
assign pbo = ~PBO;  //complement 
assign BBG = ~bbg;  //complement 
assign BBO = ~bbo;  //complement 
assign dda = ~DDA;  //complement 
assign pcg = ~PCG;  //complement 
assign BCG = ~bcg;  //complement 
assign BCO = ~bco;  //complement 
assign ddb = ~DDB;  //complement 
assign pco = ~PCO;  //complement 
assign BDG = ~bdg;  //complement 
assign BDO = ~bdo;  //complement 
assign ddc = ~DDC;  //complement 
assign pdg = ~PDG;  //complement 
assign FDO = QTD & BDO ; 
assign fdo = ~FDO ; //complement 
assign FDG = QTD & BDG ; 
assign fdg = ~FDG ;  //complement 
assign FCO = QTC & BCO ; 
assign fco = ~FCO ; //complement 
assign ddd = ~DDD;  //complement 
assign pdo = ~PDO;  //complement 
assign JHG =  QVB & xae & xaf  ; 
assign jhg = ~JHG;  //complement  
assign qnc = ~QNC;  //complement 
assign MDA = ~mda;  //complement 
assign MDB = ~mdb;  //complement 
assign QME = ~qme;  //complement 
assign wag = ~WAG;  //complement 
assign wao = ~WAO;  //complement 
assign MDC = ~mdc;  //complement 
assign MDD = ~mdd;  //complement 
assign wbg = ~WBG;  //complement 
assign wbo = ~WBO;  //complement 
assign qmf = ~QMF;  //complement 
assign QOC = ~qoc;  //complement 
assign qod = ~QOD;  //complement 
assign HAG = ~hag;  //complement 
assign HBG = ~hbg;  //complement 
assign HCG = ~hcg;  //complement 
assign HDG = ~hdg;  //complement 
assign tka = qge; 
assign TKA = ~tka; //complement 
assign tkb = qge; 
assign TKB = ~tkb;  //complement 
assign tkc = qge; 
assign TKC = ~tkc;  //complement 
assign tkd = qge; 
assign TKD = ~tkd;  //complement 
assign TEA = QAD; 
assign tea = ~TEA; //complement 
assign TEB = QAD; 
assign teb = ~TEB;  //complement 
assign TEC = QAD; 
assign tec = ~TEC;  //complement 
assign TED = QAD; 
assign ted = ~TED;  //complement 
assign gag = ~GAG;  //complement 
assign gao = ~GAO;  //complement 
assign HAO = ~hao;  //complement 
assign HBO = ~hbo;  //complement 
assign HCO = ~hco;  //complement 
assign HDO = ~hdo;  //complement 
assign qge = ~QGE;  //complement 
assign qgf = ~QGF;  //complement 
assign qad = ~QAD;  //complement 
assign QOA = ~qoa;  //complement 
assign QOB = ~qob;  //complement 
assign gbg = ~GBG;  //complement 
assign gbo = ~GBO;  //complement 
assign tqd =  qao & qae  ; 
assign TQD = ~tqd;  //complement 
assign wcg = ~WCG;  //complement 
assign wco = ~WCO;  //complement 
assign kag = ~KAG;  //complement 
assign kao = ~KAO;  //complement 
assign wdg = ~WDG;  //complement 
assign wdo = ~WDO;  //complement 
assign JEG =  LBA & lbb & lbc & lbd & lbe & lbf  ; 
assign jeg = ~JEG;  //complement  
assign mca = ~MCA;  //complement 
assign mcb = ~MCB;  //complement 
assign mcc = ~MCC;  //complement 
assign mde = ~MDE;  //complement 
assign mba = ~MBA;  //complement 
assign mbb = ~MBB;  //complement 
assign mbc = ~MBC;  //complement 
assign OAG = ~oag;  //complement 
assign OAO = ~oao;  //complement 
assign OEG = ~oeg;  //complement 
assign QMH = ~qmh;  //complement 
assign gcg = ~GCG;  //complement 
assign gco = ~GCO;  //complement 
assign eag = ~EAG;  //complement 
assign eao = ~EAO;  //complement 
assign maa = ~MAA;  //complement 
assign mab = ~MAB;  //complement 
assign mac = ~MAC;  //complement 
assign nag = ~NAG;  //complement 
assign nao = ~NAO;  //complement 
assign lag = ~LAG;  //complement 
assign sag = ~SAG;  //complement 
assign OBG = ~obg;  //complement 
assign OBO = ~obo;  //complement 
assign OEO = ~oeo;  //complement 
assign nbg = ~NBG;  //complement 
assign nbo = ~NBO;  //complement 
assign thc =  qgd & qhd  ; 
assign THC = ~thc;  //complement 
assign AAG = ~aag;  //complement 
assign ABG = ~abg;  //complement 
assign ABO = ~abo;  //complement 
assign okg = ~OKG;  //complement 
assign ncg = ~NCG;  //complement 
assign nco = ~NCO;  //complement 
assign JJA =  QAB & cap & cao & CAN  ; 
assign jja = ~JJA;  //complement  
assign JKG =  cam & CAL & CAK & caj  ; 
assign jkg = ~JKG;  //complement 
assign AAO = ~aao;  //complement 
assign CAO = ~cao;  //complement 
assign oko = ~OKO;  //complement 
assign ndg = ~NDG;  //complement 
assign ndo = ~NDO;  //complement 
assign qga = ~QGA;  //complement 
assign qua = ~QUA;  //complement 
assign okt = ~OKT;  //complement 
assign qqb = ~QQB;  //complement 
assign OCG = ~ocg;  //complement 
assign OCO = ~oco;  //complement 
assign OFG = ~ofg;  //complement 
assign qgb = ~QGB;  //complement 
assign qgc = ~QGC;  //complement 
assign gdg = ~GDG;  //complement 
assign gdo = ~GDO;  //complement 
assign ebg = ~EBG;  //complement 
assign ebo = ~EBO;  //complement 
assign olf = ~OLF;  //complement 
assign qgd = ~QGD;  //complement 
assign ODG = ~odg;  //complement 
assign ODO = ~odo;  //complement 
assign OFO = ~ofo;  //complement 
assign VAB = ~vab;  //complement 
assign pah = ~PAH;  //complement 
assign xah = ~XAH;  //complement 
assign pap = ~PAP;  //complement 
assign FAH = QTA & BAH ; 
assign fah = ~FAH ; //complement 
assign FAP = QTA & BAP ; 
assign fap = ~FAP ;  //complement 
assign FBH = QTB & BBH ; 
assign fbh = ~FBH ;  //complement 
assign FBP = QTB & BBP; 
assign fbp = ~FBP; 
assign pdp = ~PDP;  //complement 
assign pbh = ~PBH;  //complement 
assign BAH = ~bah;  //complement 
assign BAP = ~bap;  //complement 
assign VDB = ~vdb;  //complement 
assign pbp = ~PBP;  //complement 
assign BBH = ~bbh;  //complement 
assign BBP = ~bbp;  //complement 
assign vad = ~VAD;  //complement 
assign pch = ~PCH;  //complement 
assign BCH = ~bch;  //complement 
assign BCP = ~bcp;  //complement 
assign vbd = ~VBD;  //complement 
assign pcp = ~PCP;  //complement 
assign BDH = ~bdh;  //complement 
assign BDP = ~bdp;  //complement 
assign vcd = ~VCD;  //complement 
assign VBB = ~vbb;  //complement 
assign VCB = ~vcb;  //complement 
assign pdh = ~PDH;  //complement 
assign FDP = QTD & BDP ; 
assign fdp = ~FDP ; //complement 
assign FDH = QTD & BDH ; 
assign fdh = ~FDH ;  //complement 
assign FCH = QTC & BCH ; 
assign fch = ~FCH ; //complement 
assign FCP = QTC & BCP ; 
assign fcp = ~FCP ;  //complement 
assign vdd = ~VDD;  //complement 
assign JHH =  QVB & xae & xaf & xag  ; 
assign jhh = ~JHH;  //complement  
assign JIB =  xae & xaf & xag & xah  ; 
assign jib = ~JIB;  //complement 
assign lca = ~LCA;  //complement 
assign qta = ~QTA;  //complement 
assign qtb = ~QTB;  //complement 
assign wah = ~WAH;  //complement 
assign wap = ~WAP;  //complement 
assign lcc = ~LCC;  //complement 
assign wbh = ~WBH;  //complement 
assign wbp = ~WBP;  //complement 
assign HAH = ~hah;  //complement 
assign HBH = ~hbh;  //complement 
assign HCH = ~hch;  //complement 
assign HDH = ~hdh;  //complement 
assign TMA = qge & qle ; 
assign tma = ~TMA ; //complement 
assign TMB = qge & qle ; 
assign tmb = ~TMB ;  //complement 
assign TMC = qge & qke ; 
assign tmc = ~TMC ;  //complement 
assign TMD = qge & qke; 
assign tmd = ~TMD; 
assign qke = ~QKE;  //complement 
assign qle = ~QLE;  //complement 
assign qmi = ~QMI;  //complement 
assign gah = ~GAH;  //complement 
assign gap = ~GAP;  //complement 
assign HAP = ~hap;  //complement 
assign HBP = ~hbp;  //complement 
assign HCP = ~hcp;  //complement 
assign HDP = ~hdp;  //complement 
assign tla = qld; 
assign TLA = ~tla; //complement 
assign tlb = qld; 
assign TLB = ~tlb;  //complement 
assign tlc = qkd; 
assign TLC = ~tlc;  //complement 
assign tld = qkd; 
assign TLD = ~tld;  //complement 
assign qkd = ~QKD;  //complement 
assign qld = ~QLD;  //complement 
assign gbh = ~GBH;  //complement 
assign gbp = ~GBP;  //complement 
assign wch = ~WCH;  //complement 
assign wcp = ~WCP;  //complement 
assign kah = ~KAH;  //complement 
assign kap = ~KAP;  //complement 
assign qtc = ~QTC;  //complement 
assign wdh = ~WDH;  //complement 
assign wdp = ~WDP;  //complement 
assign qkb = ~QKB;  //complement 
assign qlb = ~QLB;  //complement 
assign qlc = ~QLC;  //complement 
assign lcb = ~LCB;  //complement 
assign JGD =  QMG & lca & lcb & lcc  ; 
assign jgd = ~JGD;  //complement  
assign JGE =  lca & lcb & lcc & lcd  ; 
assign jge = ~JGE;  //complement 
assign JGC =  QMG & lca & lcb  ; 
assign jgc = ~JGC;  //complement 
assign JGA =  QMG  ; 
assign jga = ~JGA;  //complement 
assign JGB =  QMG & lca  ; 
assign jgb = ~JGB;  //complement 
assign OAH = ~oah;  //complement 
assign OAP = ~oap;  //complement 
assign OEH = ~oeh;  //complement 
assign lcd = ~LCD;  //complement 
assign gch = ~GCH;  //complement 
assign gcp = ~GCP;  //complement 
assign eah = ~EAH;  //complement 
assign eap = ~EAP;  //complement 
assign qha = ~QHA;  //complement 
assign nah = ~NAH;  //complement 
assign nap = ~NAP;  //complement 
assign lah = ~LAH;  //complement 
assign sah = ~SAH;  //complement 
assign OBH = ~obh;  //complement 
assign OBP = ~obp;  //complement 
assign OEP = ~oep;  //complement 
assign nbh = ~NBH;  //complement 
assign nbp = ~NBP;  //complement 
assign JGG =  laa & lab & lac & lad & lae & laf  ; 
assign jgg = ~JGG;  //complement  
assign AAH = ~aah;  //complement 
assign AAR = ~aar;  //complement 
assign ABH = ~abh;  //complement 
assign qab = ~QAB;  //complement 
assign okh = ~OKH;  //complement 
assign nch = ~NCH;  //complement 
assign ncp = ~NCP;  //complement 
assign JKH =  cam & CAL & CAK & CAJ  ; 
assign jkh = ~JKH;  //complement  
assign AAP = ~aap;  //complement 
assign ABP = ~abp;  //complement 
assign CAP = ~cap;  //complement 
assign okp = ~OKP;  //complement 
assign ndh = ~NDH;  //complement 
assign ndp = ~NDP;  //complement 
assign qhe = ~QHE;  //complement 
assign jma =  qat & qaa  ; 
assign JMA = ~jma;  //complement 
assign jmb =  qat & qaa  ; 
assign JMB = ~jmb;  //complement 
assign OCH = ~och;  //complement 
assign OCP = ~ocp;  //complement 
assign OFH = ~ofh;  //complement 
assign okr = ~OKR;  //complement 
assign qhb = ~QHB;  //complement 
assign qhc = ~QHC;  //complement 
assign gdh = ~GDH;  //complement 
assign gdp = ~GDP;  //complement 
assign ebh = ~EBH;  //complement 
assign ebp = ~EBP;  //complement 
assign olg = ~OLG;  //complement 
assign qhd = ~QHD;  //complement 
assign ODH = ~odh;  //complement 
assign ODP = ~odp;  //complement 
assign OFP = ~ofp;  //complement 
assign qat = ~QAT;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iff = ~IFF; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign iki = ~IKI; //complement 
assign ikj = ~IKJ; //complement 
assign ikk = ~IKK; //complement 
assign ikl = ~IKL; //complement 
assign ikm = ~IKM; //complement 
assign ikn = ~IKN; //complement 
assign iko = ~IKO; //complement 
assign ikp = ~IKP; //complement 
assign ikq = ~IKQ; //complement 
assign ikr = ~IKR; //complement 
assign iks = ~IKS; //complement 
assign ikt = ~IKT; //complement 
assign ima = ~IMA; //complement 
assign ina = ~INA; //complement 
assign inb = ~INB; //complement 
assign inc = ~INC; //complement 
assign ind = ~IND; //complement 
always@(posedge IZZ )
   begin 
 vaa <= qna ; 
 PAA <=  RAA & TAA  |  REA & TBA  |  RIA & TCA  |  RMA & TDA  |  FAA  ; 
 XAA <=  XAA & tta & jha  |  xaa & JHA  ; 
 vba <= qnb ; 
 PAI <=  RAI & TAB  |  REI & TBB  |  RII & TCB  |  RMI & TDB  |  FAI  ; 
 vca <= qnc ; 
 PBA <=  RBA & TAC  |  RFA & TBC  |  RJA & TCC  |  RNA & TDC  |  FBA  ; 
 baa <=  waa & TKA  |  haa & TLA  |  baa & TMA  ; 
 bai <=  wai & TKA  |  hai & TLA  |  bai & TMA  ; 
 vda <= qnd ; 
 PBI <=  RBI & TAD  |  RFI & TBD  |  RJI & TCD  |  RNI & TDD  |  FBI  ; 
 bba <=  wba & TKB  |  hba & TLB  |  bba & TMB  ; 
 bbi <=  wbi & TKB  |  hbi & TLB  |  bbi & TMB  ; 
 VAC <= QNA ; 
 PCA <=  RCA & TAE  |  RGA & TBE  |  RKA & TCE  |  ROA & TDE  |  FCA  ; 
 bca <=  wca & TKC  |  haa & TLC  |  bca & TMC  ; 
 bci <=  wci & TKC  |  hai & TLC  |  bci & TMC  ; 
 VBC <= QNB ; 
 PCI <=  RCI & TAF  |  RGI & TBF  |  RKI & TCF  |  ROI & TDF  |  FCI  ; 
 bda <=  wda & TKD  |  hba & TLD  |  bda & TMD  ; 
 bdi <=  wdi & TKD  |  hbi & TLD  |  bdi & TMD  ; 
 VCC <= QNC ; 
 PDA <=  RDA & TAG  |  RHA & TBG  |  RLA & TCG  |  RPA & TDG  |  FDA  ; 
 VDC <= QND ; 
 PDI <=  RDI & TAH  |  RHI & TBH  |  RLI & TCH  |  RPI & TDH  |  FDI  ; 
 LBA <=  LBA & jea & tif  |  JEA & lba  |  JFA & TIF  ; 
 LBI <=  LBA & jea & tif  |  JEA & lba  |  JFA & TIF  ; 
 WAA <=  IAA & TEA  |  HAA & TFA  ; 
 WAI <=  IAE & TEA  |  HAI & TFA  ; 
 WBA <=  IBA & TEB  |  HBA & TFB  ; 
 WBI <=  IBI & TEB  |  HBI & TFB  ; 
 haa <= aaa ; 
 hba <= haa ; 
 hca <= hba ; 
 hda <= hca ; 
 qaq <= qcj ; 
 QQE <= QDH ; 
 QTD <= JOA ; 
 QAJ <=  JQB & QAI  ; 
 QRG <=  QRF & QAI  ; 
 GAA <=  GAA & TPA  |  AAA & TPC  |  GAB & TPE  ; 
 GAI <=  GAI & TPA  |  AAI & TPC  |  GAJ & TPE  ; 
 hai <= aai ; 
 hbi <= hai ; 
 hci <= hbi ; 
 hdi <= hci ; 
 QDD <=  QDD & qac & jma  |  QDC  |  QDO  ; 
 GBA <=  GBA & TPB  |  ABA & TPD  |  GBB & TPF  ; 
 GBI <=  GBI & TPB  |  ABI & TPD  |  GBJ & TPF  ; 
 WCA <=  ICA & TEC  |  HCA & TFC  ; 
 WCI <=  ICI & TEC  |  HCI & TFC  ; 
 KAA <=  KAA & toa  |  ABA & TOA  ; 
 KAI <=  KAI & toa  |  ABI & TOA  ; 
 QPA <=  QPA & tqc  |  QPD & TQA  |  TQB  ; 
 QPE <=  QPA & tqc  |  QPD & TQA  |  TQB  ; 
 WDA <=  IDA & TED  |  HDA & TFD  ; 
 WDI <=  IDI & TED  |  HDI & TFD  ; 
 QRE <= QRD ; 
 QRF <= QRE ; 
 QRH <= QRG ; 
 QRI <= QRH ; 
 QRJ <= QRI ; 
 QRK <= QRJ ; 
 QRL <= QRK ; 
 QRM <= QRL ; 
 oaa <= paa ; 
 oai <= pai ; 
 oea <= gca ; 
 GCA <=  GCA & tpg  |  GAA & TPG  ; 
 GCI <=  GCI & tpg  |  GAI & TPG  ; 
 EAA <=  EAA & tna  |  IEA & TNA  ; 
 EAI <=  EAI & tna  |  IEI & TNA  ; 
 OGA <=  LBI  |  THC  ; 
 NAA <=  PAA & TJA  |  PBA & TJB  |  PCA & TJC  ; 
 NAI <=  PAI & TJA  |  PBI & TJB  |  PCI & TJC  ; 
 LAI <=  LAI & tie  |  AAI & TIE  ; 
 SAA <=  SAA & TSA  |  IGA & TSC  ; 
 SAI <=  SAI & TSA  |  QAK & TSC  ; 
 oba <= pba ; 
 obi <= pbi ; 
 oei <= gci ; 
 NBA <=  PDA & TJD  |  BAA & TJE  |  BBA & TJF  ; 
 NBI <=  PDI & TJD  |  BAI & TJE  |  BBI & TJF  ; 
 qak <=  iia  |  SAI  |  SAJ  ; 
 qal <=  iib  |  SAJ  ; 
 aaa <= ika ; 
 aba <= aaa ; 
 abi <= aai ; 
 OKA <=  IKA & THA  |  NAA  |  NBA  |  NCA  |  NDA  ; 
 NCA <=  BCA & TJG  |  BDA & TJH  |  SAA & TJI  ; 
 NCI <=  BCE & TJG  |  BDI & TJH  |  SAI & TJI  ; 
 aai <= iki ; 
 qaa <= ikq ; 
 OKI <=  IKI & THB  |  NAI  |  NBI  |  NCI  |  NDI  ; 
 NDA <=  EAA & TJJ  |  EBA & TJK  |  KAA & TJL  ; 
 NDI <=  EAI & TJJ  |  EBI & TJK  |  KAI & TJL  ; 
 QAN <=  QAP & IKQ  |  QAM  ; 
 QAG <=  IIA & sai & saj  |  IIB & saj  ; 
 oca <= pca ; 
 oci <= pci ; 
 ofa <= gda ; 
 okq <= ikq ; 
 QAP <=  SAI & SAK  |  SAJ & SAL  ; 
 GDA <=  GDA & tpi  |  GBA & TPI  ; 
 GDI <=  GDI & tpi  |  GBI & TPI  ; 
 EBA <=  EBA & tnb  |  IFA & TNB  ; 
 EBI <=  EBI & tnb  |  IFI & TNB  ; 
 OKS <=  jla & IKS  |  QAQ  |  QDN  ; 
 QAC <=  IKS & IKS  ; 
 QRN <= QRM ; 
 QRO <= QRN ; 
 QRP <= QRO ; 
 QSA <= QRP ; 
 LAA <=  LAA & tie  |  AAA & TIE  ; 
 oda <= pda ; 
 odi <= pdi ; 
 ofi <= gdi ; 
 PAB <=  RAB & TAA  |  REB & TBA  |  RIB & TCA  |  RMB & TDA  |  FAB  ; 
 XAB <=  XAB & tta & jhb  |  xab & JHB  ; 
 QMA <=  QPE & TQD  |  MDA  ; 
 PAJ <=  RAJ & TAB  |  REJ & TBB  |  RIJ & TCB  |  RMJ & TDB  |  FAJ  ; 
 PBB <=  RBB & TAC  |  RFB & TBC  |  RJB & TCC  |  RNB & TDC  |  FBB  ; 
 bab <=  wab & TKA  |  hab & TLA  |  bab & TMA  ; 
 baj <=  waj & TKA  |  haj & TLA  |  baj & TMA  ; 
 PBJ <=  RBJ & TAD  |  RFJ & TBD  |  RJJ & TCD  |  RNJ & TDD  |  FBJ  ; 
 bbb <=  wbb & TKB  |  hbb & TLB  |  bbb & TMB  ; 
 bbj <=  wbj & TKB  |  hbj & TLB  |  bbj & TMB  ; 
 DAA <=  DAA & jaa & tia  |  daa & JAA  ; 
 PCB <=  RCB & TAE  |  RGB & TBE  |  RKB & TCE  |  ROB & TDE  |  FCB  ; 
 bcb <=  wcb & TKC  |  hab & TLC  |  bcb & TMC  ; 
 bcj <=  wcj & TKC  |  haj & TLC  |  bcj & TMC  ; 
 DAB <=  DAB & jab & tia  |  dab & JAB  ; 
 PCJ <=  RCJ & TAF  |  RGJ & TBF  |  RKJ & TCF  |  ROJ & TDF  |  FCJ  ; 
 bdb <=  wdb & TKD  |  hbb & TLD  |  bdb & TMD  ; 
 bdj <=  wdj & TKD  |  hbj & TLD  |  bdj & TMD  ; 
 DAC <=  DAC & jac & tia  |  dac & JAC  ; 
 PDB <=  RDB & TAG  |  RHB & TBG  |  RLB & TCG  |  RPB & TDG  |  FDB  ; 
 DAD <=  DAD & jad & tia  |  dad & JAD  ; 
 PDJ <=  RDJ & TAH  |  RHJ & TBH  |  RLJ & TCH  |  RPJ & TDH  |  FDJ  ; 
 LBB <=  LBB & jeb & tif  |  JEB & lbb  |  JFB & TIF  ; 
 LBJ <=  LBB & jeb & tif  |  JEB & lbb  |  JFB & TIF  ; 
 WAB <=  IAB & TEA  |  HAB & TFA  ; 
 WAJ <=  IAJ & TEA  |  HAJ & TFA  ; 
 WBB <=  IBB & TEB  |  HBB & TFB  ; 
 WBJ <=  IBJ & TEB  |  HBJ & TFB  ; 
 hab <= aab ; 
 hbb <= hab ; 
 hcb <= hbb ; 
 hdb <= hcb ; 
 GAB <=  GAB & TPA  |  AAB & TPC  |  GAC & TPE  ; 
 GAJ <=  GAJ & TPA  |  AAJ & TPC  |  GAK & TPE  ; 
 haj <= aaj ; 
 hbj <= haj ; 
 hcj <= hbj ; 
 hdj <= hcj ; 
 QCE <=  QCE & qmh & jma  |  QCC  |  QCT  ; 
 GBB <=  GBB & TPB  |  ABB & TPD  |  GBC & TPF  ; 
 GBJ <=  GBJ & TPB  |  ABJ & TPD  |  GBK & TPF  ; 
 WCB <=  ICB & TEC  |  HCB & TFC  ; 
 WCJ <=  ICJ & TEC  |  HCJ & TFC  ; 
 KAB <=  KAB & toa  |  ABB & TOA  ; 
 KAJ <=  KAJ & toa  |  ABJ & TOA  ; 
 QPB <=  QPB & tqc & tqb  |  QPA & TQA  ; 
 QPF <=  QPB & tqc & tqb  |  QPA & TQA  ; 
 WDB <=  IDB & TED  |  HDB & TFD  ; 
 WDJ <=  IDJ & TED  |  HDJ & TFD  ; 
 QSB <= QSA ; 
 QSC <= QSB ; 
 QSD <= QSC ; 
 QSE <= QSD ; 
 QSF <= QSE ; 
 QSG <= QSF ; 
 QSH <= QSG ; 
 QSI <= QSH ; 
 oab <= pab ; 
 oaj <= paj ; 
 oeb <= gcb ; 
 GCB <=  GCB & tpg  |  GAB & TPG  ; 
 GCJ <=  GCJ & tpg  |  GAJ & TPG  ; 
 EAB <=  EAB & tna  |  IEB & TNA  ; 
 EAJ <=  EAJ & tna  |  IEJ & TNA  ; 
 ogb <=  lbj  |  THC  ; 
 NAB <=  PAB & TJA  |  PBB & TJB  |  PCB & TJC  ; 
 NAJ <=  PAJ & TJA  |  PBJ & TJB  |  PCJ & TJC  ; 
 SAB <=  SAB & TSA  |  IGB & TSC  ; 
 SAJ <=  SAJ & TSA  |  QAL & TSC  ; 
 obb <= pbb ; 
 obj <= pbj ; 
 oej <= gcj ; 
 olb <= qce ; 
 NBB <=  PDB & TJD  |  BAB & TJE  |  BBB & TJF  ; 
 NBJ <=  PDJ & TJD  |  BAJ & TJE  |  BBJ & TJF  ; 
 aab <= ikb ; 
 abb <= aab ; 
 abj <= aaj ; 
 OKB <=  IKB & THA  |  NAB  |  NBB  |  NCB  |  NDB  ; 
 NCB <=  BCB & TJG  |  BDB & TJH  |  SAB & TJI  ; 
 NCJ <=  BCJ & TJG  |  BDJ & TJH  |  SAJ & TJI  ; 
 aaj <=  ikj  ; 
 caj <=  ikj  ; 
 cbj <=  ikj  ; 
 OKJ <=  IKJ & THB  |  NAJ  |  NBJ  |  NCJ  |  NDJ  ; 
 NDB <=  EAB & TJJ  |  EBB & TJK  |  KAB & TJL  ; 
 NDJ <=  EAJ & TJJ  |  EBJ & TJK  |  KAJ & TJL  ; 
 QIA <=  JKI & JJA  ; 
 QBA <=  JKB & JKA  ; 
 ocb <= pcb ; 
 ocj <= pcj ; 
 ofb <= gdb ; 
 old <= qdd ; 
 QBB <= QBA ; 
 QIB <= QIA ; 
 GDB <=  GDB & tpi  |  GBB & TPI  ; 
 GDJ <=  GDJ & tpi  |  GBJ & TPI  ; 
 EBB <=  EBB & tnb  |  IFB & TNB  ; 
 EBJ <=  EBJ & tnb  |  IFJ & TNB  ; 
 QSJ <= QSI ; 
 QSK <= QSJ ; 
 QSL <= QSK ; 
 QSM <= QSL ; 
 LAB <=  LAB & tie  |  AAB & TIE  ; 
 LAJ <=  LAJ & tie  |  AAJ & TIE  ; 
 odb <= pdb ; 
 odj <= pdj ; 
 ofj <= gdj ; 
 PAC <=  RAC & TAA  |  REC & TBA  |  RIC & TCA  |  RMC & TDA  |  FAC  ; 
 XAC <=  XAC & tta & jhc  |  xac & JHC  ; 
 QMB <=  QPF & TQD  |  MDB  ; 
 PAK <=  RAK & TAB  |  REK & TBB  |  RIK & TCB  |  RMK & TDB  |  FAK  ; 
 PBC <=  RBC & TAC  |  RFC & TBC  |  RJC & TCC  |  RNC & TDC  |  FBC  ; 
 bac <=  wac & TKA  |  hac & TLA  |  bac & TMA  ; 
 bak <=  wak & TKA  |  hak & TLA  |  bak & TMA  ; 
 PBK <=  RBK & TAD  |  RFK & TBD  |  RJK & TCD  |  RNK & TDD  |  FBK  ; 
 bbc <=  wbc & TKB  |  hbc & TLB  |  bbc & TMB  ; 
 bbk <=  wbk & TKB  |  hbk & TLB  |  bbk & TMB  ; 
 DBA <=  DBA & jba & tib  |  dba & JBA  ; 
 PCC <=  RCC & TAE  |  RGC & TBE  |  RKC & TCE  |  ROC & TDE  |  FCC  ; 
 bcc <=  wcc & TKC  |  hac & TLC  |  bcc & TMC  ; 
 bck <=  wck & TKC  |  hak & TLC  |  bck & TMC  ; 
 DBB <=  DBB & jbb & tib  |  dbb & JBB  ; 
 PCK <=  RCK & TAF  |  RGK & TBF  |  RKK & TCF  |  ROK & TDF  |  FCK  ; 
 bdc <=  wdc & TKD  |  hbc & TLD  |  bdc & TMD  ; 
 bdk <=  wdk & TKD  |  hbk & TLD  |  bdk & TMD  ; 
 DBC <=  DBC & jbc & tib  |  dbc & JBC  ; 
 PDC <=  RDC & TAG  |  RHC & TBG  |  RLC & TCG  |  RPC & TDG  |  FDC  ; 
 DBD <=  DBD & jbd & tib  |  dbd & JBD  ; 
 PDK <=  RDK & TAH  |  RHK & TBH  |  RLK & TCH  |  RPK & TDH  |  FDK  ; 
 QND <=  QPH & QDH  |  MDD  ; 
 LBC <=  LBC & jec & tif  |  JEC & lbc  |  JFC & TIF  ; 
 LBK <=  LBC & jec & tif  |  JEC & lbc  |  JFC & TIF  ; 
 QCG <= QCF ; 
 QCH <= QCG ; 
 QCI <= QCH ; 
 WAC <=  IAC & TEA  |  HAC & TFA  ; 
 WAK <=  IAK & TEA  |  HAK & TFA  ; 
 QCT <=  qmj & QCS  ; 
 QCU <=  QMJ & QCS  ; 
 WBC <=  IBC & TEB  |  HBC & TFB  ; 
 WBK <=  IBK & TEB  |  HBK & TFB  ; 
 QCN <= QCM ; 
 QCQ <= QCP ; 
 QCR <= QCQ ; 
 QCS <= QCR ; 
 hac <= aac ; 
 hbc <= hac ; 
 hcc <= hbc ; 
 hdc <= hcc ; 
 QCB <=  QCA & QMH  ; 
 QCF <=  QCE & QMH  ; 
 QCC <= QCB ; 
 QCJ <= QCI ; 
 QCL <= QCK ; 
 QCM <= QCL ; 
 GAC <=  GAC & TPA  |  AAC & TPC  |  GAD & TPE  ; 
 GAK <=  GAK & TPA  |  AAK & TPC  |  GAL & TPE  ; 
 hak <= aak ; 
 hbk <= hak ; 
 hck <= hbk ; 
 hdk <= hck ; 
 QCO <=  QCO & gac & jma  |  QCN & JEG  ; 
 QCK <=  QCJ & QAC  |  QCN & jeg  ; 
 QCP <=  QCO & QAC  ; 
 GBC <=  GBC & TPB  |  ABC & TPD  |  GBD & TPF  ; 
 GBK <=  GBK & TPB  |  ABK & TPD  |  GBL & TPF  ; 
 WCC <=  ICC & TEC  |  HCC & TFC  ; 
 WCK <=  ICK & TEC  |  HCK & TFC  ; 
 KAC <=  KAC & toa  |  ABC & TOA  ; 
 KAK <=  KAK & toa  |  ABK & TOA  ; 
 QPC <=  QPC & tqc & tqb  |  QPB & TQA  ; 
 QPG <=  QPC & tqc & tqb  |  QPB & TQA  ; 
 WDC <=  IDC & TED  |  HDC & TFD  ; 
 WDK <=  IDK & TED  |  HDK & TFD  ; 
 QKC <= QKB ; 
 oac <= pac ; 
 oak <= pak ; 
 oec <= gcc ; 
 GCC <=  GCC & tpg  |  GAC & TPG  ; 
 GCK <=  GCK & tpg  |  GAK & TPG  ; 
 EAC <=  EAC & tna  |  IEC & TNA  ; 
 EAK <=  EAK & tna  |  IEK & TNA  ; 
 ogc <=  lbk  |  THC  ; 
 NAC <=  PAC & TJA  |  PBC & TJB  |  PCC & TJC  ; 
 NAK <=  PAK & TJA  |  PBK & TJB  |  PCK & TJC  ; 
 LAC <=  LAC & tie  |  AAC & TIE  ; 
 SAC <=  SAC & TSA  |  IGC & TSC  ; 
 obc <= pbc ; 
 obk <= pbk ; 
 oek <= gck ; 
 QJB <= QJA ; 
 NBC <=  PDC & TJD  |  BAC & TJE  |  BBC & TJF  ; 
 NBK <=  PDK & TJD  |  BAK & TJE  |  BBK & TJF  ; 
 aac <= ikc ; 
 abc <= aac ; 
 abk <= aak ; 
 OKC <=  IKC & THA  |  NAC  |  NBC  |  NCC  |  NDC  ; 
 NCC <=  BCC & TJG  |  BDC & TJH  |  SAC & TJI  ; 
 NCK <=  BCK & TJG  |  BDK & TJH  |  SAK & TJI  ; 
 aak <=  ikk  ; 
 cak <=  ikk  ; 
 cbk <=  ikk  ; 
 OKK <=  IKK & THB  |  NAK  |  NBK  |  NCK  |  NDK  ; 
 NDC <=  EAC & TJJ  |  EBC & TJK  |  KAC & TJL  ; 
 NDK <=  EAK & TJJ  |  EBK & TJK  |  KAK & TJL  ; 
 QCA <=  JKC & JJA  ; 
 QJA <=  JKJ & JJA  ; 
 SAK <=  SAK & tsb  |  ABA & TSB  ; 
 occ <= pcc ; 
 ock <= pck ; 
 ofc <= gdc ; 
 olc <= qco ; 
 GDC <=  GDC & tpi  |  GBC & TPI  ; 
 GDK <=  GDK & tpi  |  GBK & TPI  ; 
 EBC <=  EBC & tnb  |  IFC & TNB  ; 
 EBK <=  EBK & tnb  |  IFK & TNB  ; 
 odc <= pdc ; 
 odk <= pdk ; 
 ofk <= gdk ; 
 uaa <= daa ; 
 uab <= dab ; 
 uac <= dac ; 
 uad <= dad ; 
 PAD <=  RAD & TAA  |  RED & TBA  |  RID & TCA  |  RMD & TDA  |  FAD  ; 
 XAD <=  XAD & tta & jhd  |  xad & JHD  ; 
 uai <= daa ; 
 uaj <= dab ; 
 uak <= dac ; 
 ual <= dad ; 
 PAL <=  RAL & TAB  |  REL & TBB  |  RIL & TCB  |  RML & TDB  |  FAL  ; 
 uba <= dba ; 
 ubb <= dbb ; 
 ubc <= dbc ; 
 ubd <= dbd ; 
 PBD <=  RBD & TAC  |  RFD & TBC  |  RJD & TCC  |  RND & TDC  |  FBD  ; 
 bad <=  wad & TKA  |  had & TLA  |  bad & TMA  ; 
 bal <=  wal & TKA  |  hal & TLA  |  bal & TMA  ; 
 ubi <= dba ; 
 ubj <= dbb ; 
 ubk <= dbc ; 
 ubl <= dbd ; 
 PBL <=  RBL & TAD  |  RFL & TBD  |  RJL & TCD  |  RNL & TDD  |  FBL  ; 
 bbd <=  wbd & TKB  |  hbd & TLB  |  bbd & TMB  ; 
 bbl <=  wbl & TKB  |  hbl & TLB  |  bbl & TMB  ; 
 uca <= dca ; 
 ucb <= dcb ; 
 ucc <= dcc ; 
 ucd <= dcd ; 
 PCD <=  RCD & TAE  |  RGD & TBE  |  RKD & TCE  |  ROD & TDE  |  FCD  ; 
 bcd <=  wcd & TKC  |  had & TLC  |  bcd & TMC  ; 
 bcl <=  wcl & TKC  |  hal & TLC  |  bcl & TMC  ; 
 uci <= dca ; 
 ucj <= dcb ; 
 uck <= dcc ; 
 ucl <= dcd ; 
 PCL <=  RCL & TAF  |  RGL & TBF  |  RKL & TCF  |  ROL & TDF  |  FCL  ; 
 bdd <=  wdd & TKD  |  hbd & TLD  |  bdd & TMD  ; 
 bdl <=  wdl & TKD  |  hbl & TLD  |  bdl & TMD  ; 
 uda <= dda ; 
 udb <= ddb ; 
 udc <= ddc ; 
 udd <= ddd ; 
 PDD <=  RDD & TAG  |  RHD & TBG  |  RLD & TCG  |  RPD & TDG  |  FDD  ; 
 udi <= dda ; 
 udj <= ddb ; 
 udk <= ddc ; 
 udl <= ddd ; 
 PDL <=  RDL & TAH  |  RHL & TBH  |  RLL & TCH  |  RPL & TDH  |  FDL  ; 
 LBD <=  LBD & jed & tif  |  JED & lbd  |  JFD & TIF  ; 
 LBL <=  LBD & jed & tif  |  JED & lbd  |  JFD & TIF  ; 
 WAD <=  IAD & TEA  |  HAD & TFA  ; 
 WAL <=  IAL & TEA  |  HAL & TFA  ; 
 QDB <= QDA ; 
 QDC <= QDB ; 
 QDF <= QDE ; 
 QDG <= QDF ; 
 WBD <=  IBD & TEB  |  HBD & TFB  ; 
 WBL <=  IBL & TEB  |  HBL & TFB  ; 
 QDH <= QDG ; 
 QDL <= QDK ; 
 QDM <= QDL ; 
 QDN <= QDM ; 
 had <= aad ; 
 hbd <= had ; 
 hcd <= hbd ; 
 hdd <= hcd ; 
 QDO <=  QDN & qmj  ; 
 QDE <=  QDD & QAC  |  qmf & QDH  ; 
 GAD <=  GAD & TPA  |  AAD & TPC  |  GAE & TPE  ; 
 GAL <=  GAL & TPA  |  AAL & TPC  |  GAM & TPE  ; 
 hal <= aal ; 
 hbl <= hal ; 
 hcl <= hbl ; 
 hdl <= hcl ; 
 QDJ <=  QDJ & qaf & jma  |  QDI  ; 
 QDK <=  QDJ & QAF  ; 
 QMG <=  QCP & QAF  |  QDK  ; 
 GBD <=  GBD & TPB  |  ABD & TPD  |  GBE & TPF  ; 
 GBL <=  GBL & TPB  |  ABL & TPD  |  GBM & TPF  ; 
 QDI <= QDH & QMF ; 
 WCD <=  ICD & TEC  |  HCD & TFC  ; 
 WCL <=  ICL & TEC  |  HCL & TFC  ; 
 KAD <=  KAD & toa  |  ABD & TOA  ; 
 KAL <=  KAL & toa  |  ABL & TOA  ; 
 QPD <=  QPD & tqc & tqb  |  QPC & TQA  ; 
 QPH <=  QPD & tqc & tqb  |  QPC & TQA  ; 
 WDD <=  IDD & TED  |  HDD & TFD  ; 
 WDL <=  IDL & TED  |  HDL & TFD  ; 
 QRA <= QAH ; 
 QRB <= QRA ; 
 QRC <= QRB ; 
 QRD <= QRC ; 
 QSN <= QSM ; 
 QSO <= QSN ; 
 QSP <= QSO ; 
 oge <=  lbm  |  THC  ; 
 oad <= pad ; 
 oal <= pal ; 
 oed <= gcd ; 
 GCD <=  GCD & tpg  |  GAD & TPG  ; 
 GCL <=  GCL & tpg  |  GAL & TPG  ; 
 EAD <=  EAD & tna  |  IED & TNA  ; 
 EAL <=  EAL & tna  |  IEL & TNA  ; 
 ogd <=  lbl  |  THC  ; 
 OHB <=  QCC  |  QCT  |  QGC  ; 
 NAD <=  PAD & TJA  |  PBD & TJB  |  PCD & TJC  ; 
 NAL <=  PAL & TJA  |  PBL & TJB  |  PCL & TJC  ; 
 LAD <=  LAD & tie  |  AAD & TIE  ; 
 SAD <=  SAD & TSA  |  IGD & TSC  ; 
 obd <= pbd ; 
 obl <= pbl ; 
 oel <= gcl ; 
 NBD <=  PDD & TJD  |  BAD & TJE  |  BBD & TJF  ; 
 NBL <=  PDL & TJD  |  BAL & TJE  |  BBL & TJF  ; 
 OHA <=  QCC  |  QCT  |  QDI  |  QGC  |  JLD  ; 
 QAH <=  QCC  |  QCT  |  QDI  |  QGC  |  JLD  ; 
 aad <= ikd ; 
 abd <= aad ; 
 abl <= aal ; 
 ole <= qdj ; 
 OKD <=  IKD & THA  |  NAD  |  NBD  |  NCD  |  NDD  ; 
 NCD <=  BCD & TJG  |  BDD & TJH  |  SAD & TJI  ; 
 NCL <=  BCL & TJG  |  BDL & TJH  |  SAL & TJI  ; 
 aal <=  ikl  ; 
 cal <=  ikl  ; 
 cbl <=  ikl  ; 
 OKL <=  IKL & THB  |  NAL  |  NBL  |  NCL  |  NDL  ; 
 NDD <=  EAD & TJJ  |  EBD & TJK  |  KAD & TJL  ; 
 NDL <=  EAL & TJJ  |  EBL & TJK  |  KAL & TJL  ; 
 QDA <=  JKD & JJA  ; 
 QKA <=  JKK & JJA  ; 
 SAL <=  SAL & tsb  |  ABB & TSB  ; 
 ocd <= pcd ; 
 ocl <= pcl ; 
 ofd <= gdd ; 
 QAF <= IJB ; 
 GDD <=  GDD & tpi  |  GBD & TPI  ; 
 GDL <=  GDL & tpi  |  GBL & TPI  ; 
 EBD <=  EBD & tnb  |  IFD & TNB  ; 
 EBL <=  EBL & tnb  |  IFL & TNB  ; 
 OLA <=  QAI & qsp & jmb  |  QAH  ; 
 QAI <=  QAI & qsp & jmb  |  QAH  ; 
 odd <= pdd ; 
 odl <= pdl ; 
 ofl <= gdl ; 
 uae <= daa ; 
 uaf <= dab ; 
 uag <= dac ; 
 uah <= dad ; 
 PAE <=  RAE & TAA  |  REE & TBA  |  RIE & TCA  |  RME & TDA  |  FAE  ; 
 XAE <=  XAE & tta & jhe  |  xae & JHE  ; 
 uam <= daa ; 
 uan <= dab ; 
 uao <= dac ; 
 uap <= dad ; 
 PAM <=  RAM & TAB  |  REM & TBB  |  RIM & TCB  |  RMM & TDB  |  FAM  ; 
 ube <= dba ; 
 ubf <= dbb ; 
 ubg <= dbc ; 
 ubh <= dbd ; 
 PBE <=  RBE & TAC  |  RFE & TBC  |  RJE & TCC  |  RNE & TDC  |  FBE  ; 
 bae <=  wae & TKA  |  hae & TLA  |  bae & TMA  ; 
 bam <=  wam & TKA  |  ham & TLA  |  bam & TMA  ; 
 ubm <= dba ; 
 ubn <= dbb ; 
 ubo <= dbc ; 
 ubp <= dbd ; 
 PBM <=  RBM & TAD  |  RFM & TBD  |  RJM & TCD  |  RNM & TDD  |  FBM  ; 
 bbe <=  wbe & TKB  |  hbe & TLB  |  bbe & TMB  ; 
 bbm <=  wbm & TKB  |  hbm & TLB  |  bbm & TMB  ; 
 uce <= dca ; 
 ucf <= dcb ; 
 ucg <= dcc ; 
 uch <= dcd ; 
 PCE <=  RCE & TAE  |  RGE & TBE  |  RKE & TCE  |  ROE & TDE  |  FCE  ; 
 bce <=  wce & TKC  |  hae & TLC  |  bce & TMC  ; 
 bcm <=  wcm & TKC  |  ham & TLC  |  bcm & TMC  ; 
 ucm <= dca ; 
 ucn <= dcb ; 
 uco <= dcc ; 
 ucp <= dcd ; 
 PCM <=  RCM & TAF  |  RGM & TBF  |  RKM & TCF  |  ROM & TDF  |  FCM  ; 
 bde <=  wde & TKD  |  hbe & TLD  |  bde & TMD  ; 
 bdm <=  wdm & TKD  |  hbm & TLD  |  bdm & TMD  ; 
 ude <= dda ; 
 udf <= ddb ; 
 udg <= ddc ; 
 udh <= ddd ; 
 WDE <=  IDE & TED  |  HDE & TFD  ; 
 udm <= dda ; 
 udn <= ddb ; 
 udo <= ddc ; 
 udp <= ddd ; 
 PDM <=  RDM & TAH  |  RHM & TBH  |  RLM & TCH  |  RPM & TDH  |  FDM  ; 
 QNA <=  QPE & QDH  |  MDA  ; 
 LBE <=  LBE & jee & tif  |  JEE & lbe  |  JFE & TIF  ; 
 LBM <=  LBE & jee & tif  |  JEE & lbe  |  JFE & TIF  ; 
 WAE <=  IAE & TEA  |  HAE & TFA  ; 
 WAM <=  IAM & TEA  |  HAM & TFA  ; 
 QQA <=  JLB  |  JLC  |  QUC  ; 
 WBE <=  IBE & TEB  |  HBE & TFB  ; 
 WBM <=  IBM & TEB  |  HBM & TFB  ; 
 hae <= aae ; 
 hbe <= hae ; 
 hce <= hbe ; 
 hde <= hce ; 
 GAE <=  GAE & TPA  |  AAE & TPC  |  GAF & TPE  ; 
 GAM <=  GAM & TPA  |  AAM & TPC  |  GAN & TPE  ; 
 ham <= aam ; 
 hbm <= ham ; 
 hcm <= hbm ; 
 hdm <= hcm ; 
 QQD <=  QQD & qqc & jma  |  QOA  ; 
 QAE <= IJA ; 
 QQC <= QQB ; 
 GBE <=  GBE & TPB  |  ABE & TPD  |  GBF & TPF  ; 
 GBM <=  GBM & TPB  |  ABM & TPD  |  GBN & TPF  ; 
 WCE <=  ICE & TEC  |  HCE & TFC  ; 
 WCM <=  ICM & TEC  |  HCM & TFC  ; 
 KAE <=  KAE & toa  |  ABE & TOA  ; 
 KAM <=  KAM & toa  |  ABM & TOA  ; 
 QMJ <=  QMI  |  JGE & JGG  ; 
 QAO <= JOB ; 
 WDM <=  IDM & TED  |  HDM & TFD  ; 
 PDE <=  RDE & TAG  |  RHE & TBG  |  RLE & TCG  |  RPE & TDG  |  FDE  ; 
 oae <= pae ; 
 oam <= pam ; 
 oee <= gce ; 
 EAE <=  EAE & tna  |  IEE & TNA  ; 
 EAM <=  EAM & tna  |  IEM & TNA  ; 
 NAE <=  PAE & TJA  |  PBE & TJB  |  PCE & TJC  ; 
 NAM <=  PAM & TJA  |  PBM & TJB  |  PCM & TJC  ; 
 LAE <=  LAE & tie  |  AAE & TIE  ; 
 SAE <=  SAE & TSA  |  IGE & TSC  ; 
 obe <= pbe ; 
 obm <= pbm ; 
 oem <= gcm ; 
 OHG <= ZZI ; 
 NBE <=  PDE & TJD  |  BAE & TJE  |  BBE & TJF  ; 
 NBM <=  PDM & TJD  |  BAM & TJE  |  BBM & TJF  ; 
 aae <= ike ; 
 abe <= aae ; 
 abm <= aam ; 
 OKE <=  IKE & THA  |  NAE  |  NBE  |  NCE  |  NDE  ; 
 NCE <=  BCE & TJG  |  BDE & TJH  |  SAE & TJI  ; 
 NCM <=  BCM & TJG  |  BDM & TJH  ; 
 aam <=  ikm  ; 
 cam <=  ikm  ; 
 cbm <=  ikm  ; 
 OKM <=  IKM & THB  |  NAM  |  NBM  |  NCM  |  NDM  ; 
 NDE <=  EAE & TJJ  |  EBE & TJK  |  KAE & TJL  ; 
 NDM <=  EAM & TJJ  |  EBM & TJK  |  KAM & TJL  ; 
 QEA <=  JKE & JJA  ; 
 QLA <=  JKL & JJA  ; 
 oce <= pce ; 
 ocm <= pcm ; 
 ofe <= gde ; 
 QEB <= QEA ; 
 GDE <=  GDE & tph  |  GBE & TPH  ; 
 GDM <=  GDM & tph  |  GBM & TPH  ; 
 EBE <=  EBE & tnb  |  IFE & TNB  ; 
 EBM <=  EBM & tnb  |  IFM & TNB  ; 
 OHD <= QUG ; 
 OHE <= QUG ; 
 OHF <= QUG ; 
 GCE <=  GCE & tpg  |  GAE & TPG  ; 
 GCM <=  GCM & tpg  |  GAM & TPG  ; 
 ode <= pde ; 
 odm <= pdm ; 
 ofm <= gdm ; 
 PAF <=  RAF & TAA  |  REF & TBA  |  RIF & TCA  |  RMF & TDA  |  FAF  ; 
 XAF <=  XAF & tta & jhf  |  xaf & JHF  ; 
 QMC <=  QPG & TQD  |  MDC  ; 
 PAN <=  RAN & TAB  |  REN & TBB  |  RIM & TCB  |  RMN & TDB  |  FAN  ; 
 PBF <=  RBF & TAC  |  RFF & TBC  |  RJF & TCC  |  RNF & TDC  |  FBF  ; 
 baf <=  waf & TKA  |  haf & TLA  |  baf & TMA  ; 
 ban <=  wan & TKA  |  han & TLA  |  ban & TMA  ; 
 PBN <=  RBN & TAD  |  RFN & TBD  |  RJN & TCD  |  RNN & TDD  |  FBN  ; 
 bbf <=  wbf & TKB  |  hbf & TLB  |  bbf & TMB  ; 
 bbn <=  wbn & TKB  |  hbn & TLB  |  bbn & TMB  ; 
 DCA <=  DCA & jca & tic  |  dca & JCA  ; 
 PCF <=  RCF & TAE  |  RGF & TBE  |  RKF & TCE  |  ROF & TDE  |  FCF  ; 
 bcf <=  wcf & TKC  |  haf & TLC  |  bcf & TMC  ; 
 bcn <=  wcn & TKC  |  han & TLC  |  bcn & TMC  ; 
 DCB <=  DCB & jcb & tic  |  dcb & JCB  ; 
 PCN <=  RCN & TAF  |  RGN & TBF  |  RKN & TCF  |  RON & TDF  |  FCN  ; 
 bdf <=  wdf & TKD  |  hbf & TLD  |  bdf & TMD  ; 
 bdn <=  wdn & TKD  |  hbn & TLD  |  bdn & TMD  ; 
 DCC <=  DCC & jcc & tic  |  dcc & JCC  ; 
 PDF <=  RDF & TAG  |  RHF & TBG  |  RLF & TCG  |  RPF & TDG  |  FDF  ; 
 DCD <=  DCD & jcd & tic  |  dcd & JCD  ; 
 PDN <=  RDN & TAH  |  RHN & TBH  |  RLN & TCH  |  RPN & TDH  |  FDN  ; 
 QNB <=  QPF & QDH  |  MDB  ; 
 LBF <=  LBF & jef & tif  |  JEF & lbf  |  JFF & TIF  ; 
 LBN <=  LBF & jef & tif  |  JEF & lbf  |  JFF & TIF  ; 
 QVB <=  QUC & JIA  ; 
 QVC <=  JIB & JIA  ; 
 WAF <=  IAF & TEA  |  HAF & TFA  ; 
 WAN <=  IAN & TEA  |  HAN & TFA  ; 
 QUB <= QUA ; 
 QVA <= QUC ; 
 WBF <=  IBF & TEB  |  HBF & TFB  ; 
 WBN <=  IBN & TEB  |  HBN & TFB  ; 
 haf <= aaf ; 
 hbf <= haf ; 
 hcf <= hbf ; 
 hdf <= hcf ; 
 QUC <=  QUB  |  QUE  ; 
 QUG <=  QUC  |  QUE  |  QUD  ; 
 GAF <=  GAF & TPA  |  AAF & TPC  |  GAG & TPE  ; 
 GAN <=  GAN & TPA  |  AAN & TPC  |  GAO & TPE  ; 
 han <= aan ; 
 hbn <= han ; 
 hcn <= hbn ; 
 hdn <= hcn ; 
 QUD <=  QUD & qaf & jma  |  QUC  ; 
 que <=  qud  |  qaf  |  QVC  ; 
 quf <=  qud  |  qaf  |  qvc  ; 
 GBF <=  GBF & TPB  |  ABF & TPD  |  GBG & TPF  ; 
 GBN <=  GBN & TPB  |  ABN & TPD  |  GBO & TPF  ; 
 QAM <=  QAP & IKQ  ; 
 WCF <=  ICF & TEC  |  HCF & TFC  ; 
 WCN <=  ICN & TEC  |  HCN & TFC  ; 
 KAF <=  KAF & toa  |  ABF & TOA  ; 
 KAN <=  KAN & toa  |  ABN & TOA  ; 
 WDF <=  IDF & TED  |  HDF & TFD  ; 
 WDN <=  IDN & TED  |  HDN & TFD  ; 
 oaf <= paf ; 
 oan <= pan ; 
 oef <= gcf ; 
 GCF <=  GCF & tpg  |  GAF & TPG  ; 
 GCN <=  GCN & tpg  |  GAN & TPG  ; 
 EAF <=  EAF & tna  |  IEF & TNA  ; 
 EAN <=  EAN & tna  |  IEN & TNA  ; 
 ogf <=  lbn  |  THC  ; 
 NAF <=  PAF & TJA  |  PBF & TJB  |  PCF & TJC  ; 
 NAN <=  PAN & TJA  |  PBN & TJB  |  PCN & TJC  ; 
 LAF <=  LAF & tie  |  AAF & TIE  ; 
 SAF <=  SAF & TSA  |  IGF & TSC  ; 
 obf <= pbf ; 
 obn <= pbn ; 
 oen <= gcn ; 
 QUH <= IND ; 
 NBF <=  PDF & TJD  |  BAF & TJE  |  BBF & TJF  ; 
 NBN <=  PDN & TJD  |  BAM & TJE  |  BBN & TJF  ; 
 OHC <=  QUG & QUH  |  INA & QUH  |  INB & QUH  |  INC & QUH  ; 
 aaf <= ikf ; 
 abf <= aaf ; 
 abn <= aan ; 
 OKF <=  IKF & THA  |  NAF  |  NBF  |  NCF  |  NDF  ; 
 NCF <=  BCF & TJG  |  BDF & TJH  |  SAF & TJI  ; 
 NCN <=  BCN & TJG  |  BDN & TJH  ; 
 aan <=  ikn  ; 
 can <=  ikn  ; 
 OKN <=  IKN & THB  |  NAN  |  NBN  |  NCN  |  NDN  ; 
 NDF <=  EAF & TJJ  |  EBF & TJK  |  KAF & TJL  ; 
 NDN <=  EAN & TJJ  |  EBN & TJK  |  KAN & TJL  ; 
 QFA <=  JJA & JKF  ; 
 QFB <=  QFA & JKF  ; 
 ocf <= pcf ; 
 ocn <= pcn ; 
 off <= gdf ; 
 olh <= qud ; 
 GDF <=  GDF & tph  |  GBF & TPH  ; 
 GDN <=  GDN & tph  |  GBN & TPH  ; 
 EBF <=  EBF & tnb  |  IFF & TNB  ; 
 EBN <=  EBN & tnb  |  IFN & TNB  ; 
 odf <= pdf ; 
 odn <= pdn ; 
 ofn <= gdn ; 
 PAG <=  RAG & TAA  |  REG & TBA  |  RIG & TCA  |  RMG & TDA  |  FAG  ; 
 XAG <=  XAG & tta & jhg  |  xag & JHG  ; 
 QMD <=  QPH & TQD  |  MDD  ; 
 PAO <=  RAO & TAB  |  REO & TBB  |  RIO & TCB  |  RMO & TDB  |  FAO  ; 
 PBG <=  RBG & TAC  |  RFG & TBC  |  RJG & TCC  |  RNG & TDC  |  FBG  ; 
 bag <=  wag & TKA  |  hag & TLA  |  bag & TMA  ; 
 bao <=  wao & TKA  |  hao & TLA  |  bao & TMA  ; 
 PBO <=  RBO & TAD  |  RFO & TBD  |  RJO & TCD  |  RNO & TDD  |  FBO  ; 
 bbg <=  wbg & TKB  |  hbg & TLB  |  bbg & TMB  ; 
 bbo <=  wbo & TKB  |  hbo & TLB  |  bbo & TMB  ; 
 DDA <=  DDA & jda & tid  |  dda & JDA  ; 
 PCG <=  RCG & TAE  |  RGG & TBE  |  RKG & TCE  |  ROG & TDE  |  FCG  ; 
 bcg <=  wcg & TKC  |  hag & TLC  |  bcg & TMC  ; 
 bco <=  wco & TKC  |  hao & TLC  |  bco & TMC  ; 
 DDB <=  DDB & jdb & tid  |  ddb & JDB  ; 
 PCO <=  RCO & TAF  |  RGO & TBF  |  RKO & TCF  |  ROO & TDF  |  FCO  ; 
 bdg <=  wdg & TKD  |  hbg & TLD  |  bdg & TMD  ; 
 bdo <=  wdo & TKD  |  hbo & TLD  |  bdo & TMD  ; 
 DDC <=  DDC & jdc & tid  |  ddc & JDC  ; 
 PDG <=  RDG & TAG  |  RHG & TBG  |  RLG & TCG  |  RPG & TDG  |  FDG  ; 
 DDD <=  DDD & jdd & tid  |  ddd & JDD  ; 
 PDO <=  RDO & TAH  |  RHO & TBH  |  RLO & TCH  |  RPO & TDH  |  FDO  ; 
 QNC <=  QPG & QDH  |  MDC  ; 
 mda <=  mcc  |  MCB  |  MCA  ; 
 mdb <=  mcc  |  MCB  |  mca  ; 
 qme <=  tqd & mde  ; 
 WAG <=  IAG & TEA  |  HAG & TFA  ; 
 WAO <=  IAO & TEA  |  HAO & TFA  ; 
 mdc <=  mcc  |  mcb  |  MCA  ; 
 mdd <=  mcc  |  mcb  |  mca  ; 
 WBG <=  IBG & TEB  |  HBG & TFB  ; 
 WBO <=  IBO & TEB  |  HBO & TFB  ; 
 QMF <= JEG ; 
 qoc <= qob ; 
 QOD <= QOB ; 
 hag <= aag ; 
 hbg <= hag ; 
 hcg <= hbg ; 
 hdg <= hcg ; 
 GAG <=  GAG & TPA  |  AAG & TPC  |  GAH & TPE  ; 
 GAO <=  GAO & TPA  |  AAO & TPC  |  GAP & TPE  ; 
 hao <= aao ; 
 hbo <= hao ; 
 hco <= hbo ; 
 hdo <= hco ; 
 QGE <=  QGD & QAD  ; 
 QGF <=  QGD & QAD  ; 
 QAD <= NDE ; 
 qoa <= jja ; 
 qob <= qoa ; 
 GBG <=  GBG & TPB  |  ABG & TPD  |  GBH & TPF  ; 
 GBO <=  GBO & TPB  |  ABO & TPD  |  GBP & TPF  ; 
 WCG <=  ICG & TEC  |  HCG & TFC  ; 
 WCO <=  ICO & TEC  |  HCO & TFC  ; 
 KAG <=  KAG & toa  |  ABG & TOA  ; 
 KAO <=  KAO & toa  |  ABO & TOA  ; 
 WDG <=  IDG & TED  |  HDG & TFD  ; 
 WDO <=  IDO & TED  |  HDO & TFD  ; 
 MCA <= MBA ; 
 MCB <= MBB ; 
 MCC <= MBC ; 
 MDE <= MCC ; 
 MBA <= MAA ; 
 MBB <= MAB ; 
 MBC <= MAC ; 
 oag <= pag ; 
 oao <= pao ; 
 oeg <= gcg ; 
 qmh <=  qme  |  jeg  ; 
 GCG <=  GCG & tpg  |  GAG & TPG  ; 
 GCO <=  GCO & tpg  |  GAO & TPG  ; 
 EAG <=  EAG & tna  |  IEG & TNA  ; 
 EAO <=  EAO & tna  |  IEO & TNA  ; 
 MAA <= IHA ; 
 MAB <= IHB ; 
 MAC <= IHC ; 
 NAG <=  PAG & TJA  |  PBG & TJB  |  PCG & TJC  ; 
 NAO <=  PAO & TJA  |  PBO & TJB  |  PCO & TJC  ; 
 LAG <=  LAG & tie  |  AAG & TIE  ; 
 SAG <=  SAG & TSA  |  IGG & TSC  ; 
 obg <= pbg ; 
 obo <= pbo ; 
 oeo <= gco ; 
 NBG <=  PDG & TJD  |  BAG & TJE  |  BBG & TJF  ; 
 NBO <=  PDO & TJD  |  BAO & TJE  |  BBO & TJF  ; 
 aag <= ikg ; 
 abg <= aag ; 
 abo <= aao ; 
 OKG <=  IKG & THA  |  NAG  |  NBG  |  NCG  |  NDG  ; 
 NCG <=  BCG & TJG  |  BDG & TJH  |  SAG & TJI  ; 
 NCO <=  BCO & TJG  |  BDO & TJH  ; 
 aao <=  iko  ; 
 cao <=  iko  ; 
 OKO <=  IKO & THB  |  NAO  |  NBO  |  NCO  |  NDO  ; 
 NDG <=  EAG & TJJ  |  EBG & TJK  |  KAG & TJL  ; 
 NDO <=  EAO & TJJ  |  EBO & TJK  |  KAO & TJL  ; 
 QGA <=  JKG & JJA  ; 
 QUA <=  JKA & JJA  ; 
 OKT <=  IKT  |  QDA  |  JNA  |  JNB  |  QUF  ; 
 QQB <=  IKT  |  QDA  |  JNA  |  JNB  |  QUF  ; 
 ocg <= pcg ; 
 oco <= pco ; 
 ofg <= gdg ; 
 QGB <= QGA ; 
 QGC <= QGB ; 
 GDG <=  GDG & tph  |  GBG & TPH  ; 
 GDO <=  GDO & tph  |  GBO & TPH  ; 
 EBG <=  EBG & tnb  |  IFG & TNB  ; 
 EBO <=  EBO & tnb  |  IFO & TNB  ; 
 OLF <=  QGD & qad & jmb  |  QGC  ; 
 QGD <=  QGD & qad & jmb  |  QGC  ; 
 odg <= pdg ; 
 odo <= pdo ; 
 ofo <= gdo ; 
 vab <= qna ; 
 PAH <=  RAH & TAA  |  REH & TBA  |  RIH & TCA  |  RMH & TDA  |  FAH  ; 
 XAH <=  XAH & tta & jhh  |  xah & JHH  ; 
 PAP <=  RAP & TAB  |  REP & TBB  |  RIP & TCB  |  RMP & TDB  |  FAP  ; 
 PDP <=  RDP & TAH  |  RHP & TBH  |  RLP & TCH  |  RPP & TDH  |  FDP  ; 
 PBH <=  RBH & TAC  |  RFH & TBC  |  RJH & TCC  |  RNH & TDC  |  FBH  ; 
 bah <=  wah & TKA  |  hah & TLA  |  bah & TMA  ; 
 bap <=  wap & TKA  |  hap & TLA  |  bap & TMA  ; 
 vdb <= qnd ; 
 PBP <=  RBP & TAD  |  RFP & TBD  |  RJP & TCD  |  RNP & TDD  |  FBP  ; 
 bbh <=  wbh & TKB  |  hbh & TLB  |  bbh & TMB  ; 
 bbp <=  wbp & TKB  |  hbp & TLB  |  bbp & TMB  ; 
 VAD <= QNA ; 
 PCH <=  RCH & TAE  |  RGH & TBE  |  RKH & TCE  |  ROH & TDE  |  FCH  ; 
 bch <=  wch & TKC  |  hah & TLC  |  bch & TMC  ; 
 bcp <=  wcp & TKC  |  hap & TLC  |  bcp & TMC  ; 
 VBD <= QNB ; 
 PCP <=  RCP & TAF  |  RGP & TBF  |  RKP & TCF  |  ROP & TDF  |  FCP  ; 
 bdh <=  wdh & TKD  |  hbh & TLD  |  bdh & TMD  ; 
 bdp <=  wdp & TKD  |  hbp & TLD  |  bdp & TMD  ; 
 VCD <= QNC ; 
 vbb <= qnb ; 
 vcb <= qnc ; 
 PDH <=  RDH & TAG  |  RHH & TBG  |  RLH & TCG  |  RPH & TDG  |  FDH  ; 
 VDD <= QND ; 
 LCA <=  LCA & jga & tig  |  JGA & lca  |  LAG & TIG  ; 
 QTA <= JOA ; 
 QTB <= JOA ; 
 WAH <=  IAH & TEA  |  HAH & TFA  ; 
 WAP <=  IAP & TEA  |  HAP & TFA  ; 
 LCC <=  LCC & jgc & tig  |  JGC & lcc  |  LAI & TIG  ; 
 WBH <=  IBH & TEB  |  HBH & TFB  ; 
 WBP <=  IBP & TEB  |  HBP & TFB  ; 
 hah <= aah ; 
 hbh <= hah ; 
 hch <= hbh ; 
 hdh <= hch ; 
 QKE <= QKC ; 
 QLE <= QLC ; 
 QMI <= JGE ; 
 GAH <=  GAH & TPA  |  AAH & TPC  |  GAI & TPE  ; 
 GAP <=  GAP & TPA  |  AAP & TPC  |  GBA & TPE  ; 
 hap <= aap ; 
 hbp <= hap ; 
 hcp <= hbp ; 
 hdp <= hcp ; 
 QKD <= QKC ; 
 QLD <= QLC ; 
 GBH <=  GBH & TPB  |  ABH & TPD  |  GBI & TPF  ; 
 GBP <=  GBP & TPB  |  ABP & TPD  |  JQA & TPF  ; 
 WCH <=  ICH & TEC  |  HCH & TFC  ; 
 WCP <=  ICP & TEC  |  HCP & TFC  ; 
 KAH <=  KAH & toa  |  ABH & TOA  ; 
 KAP <=  KAP & toa  |  ABP & TOA  ; 
 QTC <= JOA ; 
 WDH <=  IDH & TED  |  HDH & TFD  ; 
 WDP <=  IDP & TED  |  HDP & TFD  ; 
 QKB <= QKA ; 
 QLB <= QLA ; 
 QLC <= QLB ; 
 LCB <=  LCB & jgb & tig  |  JGB & lcb  |  LAH & TIG  ; 
 oah <= pah ; 
 oap <= pap ; 
 oeh <= gch ; 
 LCD <=  LCD & jgd & tig  |  JGD & lcd  |  LAJ & TIG  ; 
 GCH <=  GCH & tpg  |  GAH & TPG  ; 
 GCP <=  GCP & tpg  |  GAP & TPG  ; 
 EAH <=  EAH & tna  |  IEH & TNA  ; 
 EAP <=  EAP & tna  |  IEP & TNA  ; 
 QHA <= JKH & JJA ; 
 NAH <=  PAH & TJA  |  PBH & TJB  |  PCH & TJC  ; 
 NAP <=  PAP & TJA  |  PBP & TJB  |  PCP & TJC  ; 
 LAH <=  LAH & tie  |  AAH & TIE  ; 
 SAH <=  SAH & TSA  |  IGH & TSC  ; 
 obh <= pbh ; 
 obp <= pbp ; 
 oep <= gcp ; 
 NBH <=  PDH & TJD  |  BAH & TJE  |  BBH & TJF  ; 
 NBP <=  PDP & TJD  |  BAP & TJE  |  BBP & TJF  ; 
 aah <= ikh ; 
 aar <= ikr ; 
 abh <= aah ; 
 QAB <= AAR ; 
 OKH <=  IKH & THA  |  NAH  |  NBH  |  NCH  |  NDH  ; 
 NCH <=  BCH & TJG  |  BDH & TJH  |  SAH & TJI  ; 
 NCP <=  BCP & TJG  |  BDP & TJH  ; 
 aap <= ikp ; 
 abp <= aap ; 
 cap <= ikp ; 
 OKP <=  IKP & THB  |  NAP  |  NBP  |  NCP  |  NDP  ; 
 NDH <=  EAH & TJJ  |  EBH & TJK  |  KAH & TJL  ; 
 NDP <=  EAP & TJJ  |  EBP & TJK  |  KAP & TJL  ; 
 QHE <= QAF & QHD ; 
 och <= pch ; 
 ocp <= pcp ; 
 ofh <= gdh ; 
 OKR <= IKR ; 
 QHB <= QHA ; 
 QHC <= QHB ; 
 GDH <=  GDH & tph  |  GBH & TPH  ; 
 GDP <=  GDP & tph  |  GBP & TPH  ; 
 EBH <=  EBH & tnb  |  IFH & TNB  ; 
 EBP <=  EBP & tnb  ; 
 OLG <=  QHD & qaf & jmb  |  QHC  ; 
 QHD <=  QHD & qaf & jmb  |  QHC  ; 
 odh <= pdh ; 
 odp <= pdp ; 
 ofp <= gdp ; 
 QAT <= IMA ; 
 end 
end module
